--------------------------------------------------------------------------------
-- Entity: CartridgeROM
-- Date:2011-10-25  
-- Author: jonathansieber     
--
-- Description ${cursor}
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CartridgeROM is
	port  (
		clk : in std_logic;        -- input clock, xx MHz.
		rstn : in std_logic;
		 
        ProgramAddress : in std_logic_vector(14 downto 0);
        ProgramData : out std_logic_vector(7 downto 0);
        
        CharacterAddress : in std_logic_vector(14 downto 0);
        CharacterData : out std_logic_vector(7 downto 0)
	);
end CartridgeROM;

architecture arch of CartridgeROM is

    type prg_rom_type is array (0 to 32767) of std_logic_vector(7 downto 0);
    type chr_rom_type is array (0 to 8191) of std_logic_vector(7 downto 0);
    
    signal prg_rom : prg_rom_type;
    signal chr_rom : chr_rom_type;
begin

    process (clk) begin
        if rising_edge(clk) then
            if rstn = '0' then
                prg_rom <= (
                     0 => "01111000",
                     1 => "11011000",
                     2 => "10101001",
                     3 => "00010000",
                     4 => "10001101",
                     5 => "00000000",
                     6 => "00100000",
                     7 => "10100010",
                     8 => "11111111",
                     9 => "10011010",
                     10 => "10101101",
                     11 => "00000010",
                     12 => "00100000",
                     13 => "00010000",
                     14 => "11111011",
                     15 => "10101101",
                     16 => "00000010",
                     17 => "00100000",
                     18 => "00010000",
                     19 => "11111011",
                     20 => "10100000",
                     21 => "11111110",
                     22 => "10100010",
                     23 => "00000101",
                     24 => "10111101",
                     25 => "11010111",
                     26 => "00000111",
                     27 => "11001001",
                     28 => "00001010",
                     29 => "10110000",
                     30 => "00001100",
                     31 => "11001010",
                     32 => "00010000",
                     33 => "11110110",
                     34 => "10101101",
                     35 => "11111111",
                     36 => "00000111",
                     37 => "11001001",
                     38 => "10100101",
                     39 => "11010000",
                     40 => "00000010",
                     41 => "10100000",
                     42 => "11010110",
                     43 => "00100000",
                     44 => "11001100",
                     45 => "10010000",
                     46 => "10001101",
                     47 => "00010001",
                     48 => "01000000",
                     49 => "10001101",
                     50 => "01110000",
                     51 => "00000111",
                     52 => "10101001",
                     53 => "10100101",
                     54 => "10001101",
                     55 => "11111111",
                     56 => "00000111",
                     57 => "10001101",
                     58 => "10100111",
                     59 => "00000111",
                     60 => "10101001",
                     61 => "00001111",
                     62 => "10001101",
                     63 => "00010101",
                     64 => "01000000",
                     65 => "10101001",
                     66 => "00000110",
                     67 => "10001101",
                     68 => "00000001",
                     69 => "00100000",
                     70 => "00100000",
                     71 => "00100000",
                     72 => "10000010",
                     73 => "00100000",
                     74 => "00011001",
                     75 => "10001110",
                     76 => "11101110",
                     77 => "01110100",
                     78 => "00000111",
                     79 => "10101101",
                     80 => "01111000",
                     81 => "00000111",
                     82 => "00001001",
                     83 => "10000000",
                     84 => "00100000",
                     85 => "11101101",
                     86 => "10001110",
                     87 => "01001100",
                     88 => "01010111",
                     89 => "10000000",
                     90 => "00000001",
                     91 => "10100100",
                     92 => "11001000",
                     93 => "11101100",
                     94 => "00010000",
                     95 => "00000000",
                     96 => "01000001",
                     97 => "01000001",
                     98 => "01001100",
                     99 => "00110100",
                     100 => "00111100",
                     101 => "01000100",
                     102 => "01010100",
                     103 => "01101000",
                     104 => "01111100",
                     105 => "10101000",
                     106 => "10111111",
                     107 => "11011110",
                     108 => "11101111",
                     109 => "00000011",
                     110 => "10001100",
                     111 => "10001100",
                     112 => "10001100",
                     113 => "10001101",
                     114 => "00000011",
                     115 => "00000011",
                     116 => "00000011",
                     117 => "10001101",
                     118 => "10001101",
                     119 => "10001101",
                     120 => "10001101",
                     121 => "10001101",
                     122 => "10001101",
                     123 => "10001101",
                     124 => "10001101",
                     125 => "10001101",
                     126 => "10001101",
                     127 => "10001101",
                     128 => "00000000",
                     129 => "01000000",
                     130 => "10101101",
                     131 => "01111000",
                     132 => "00000111",
                     133 => "00101001",
                     134 => "01111111",
                     135 => "10001101",
                     136 => "01111000",
                     137 => "00000111",
                     138 => "00101001",
                     139 => "01111110",
                     140 => "10001101",
                     141 => "00000000",
                     142 => "00100000",
                     143 => "10101101",
                     144 => "01111001",
                     145 => "00000111",
                     146 => "00101001",
                     147 => "11100110",
                     148 => "10101100",
                     149 => "01110100",
                     150 => "00000111",
                     151 => "11010000",
                     152 => "00000101",
                     153 => "10101101",
                     154 => "01111001",
                     155 => "00000111",
                     156 => "00001001",
                     157 => "00011110",
                     158 => "10001101",
                     159 => "01111001",
                     160 => "00000111",
                     161 => "00101001",
                     162 => "11100111",
                     163 => "10001101",
                     164 => "00000001",
                     165 => "00100000",
                     166 => "10101110",
                     167 => "00000010",
                     168 => "00100000",
                     169 => "10101001",
                     170 => "00000000",
                     171 => "00100000",
                     172 => "11100110",
                     173 => "10001110",
                     174 => "10001101",
                     175 => "00000011",
                     176 => "00100000",
                     177 => "10101001",
                     178 => "00000010",
                     179 => "10001101",
                     180 => "00010100",
                     181 => "01000000",
                     182 => "10101110",
                     183 => "01110011",
                     184 => "00000111",
                     185 => "10111101",
                     186 => "01011010",
                     187 => "10000000",
                     188 => "10000101",
                     189 => "00000000",
                     190 => "10111101",
                     191 => "01101101",
                     192 => "10000000",
                     193 => "10000101",
                     194 => "00000001",
                     195 => "00100000",
                     196 => "11011101",
                     197 => "10001110",
                     198 => "10100000",
                     199 => "00000000",
                     200 => "10101110",
                     201 => "01110011",
                     202 => "00000111",
                     203 => "11100000",
                     204 => "00000110",
                     205 => "11010000",
                     206 => "00000001",
                     207 => "11001000",
                     208 => "10111110",
                     209 => "10000000",
                     210 => "10000000",
                     211 => "10101001",
                     212 => "00000000",
                     213 => "10011101",
                     214 => "00000000",
                     215 => "00000011",
                     216 => "10011101",
                     217 => "00000001",
                     218 => "00000011",
                     219 => "10001101",
                     220 => "01110011",
                     221 => "00000111",
                     222 => "10101101",
                     223 => "01111001",
                     224 => "00000111",
                     225 => "10001101",
                     226 => "00000001",
                     227 => "00100000",
                     228 => "00100000",
                     229 => "11010001",
                     230 => "11110010",
                     231 => "00100000",
                     232 => "01011100",
                     233 => "10001110",
                     234 => "00100000",
                     235 => "10000010",
                     236 => "10000001",
                     237 => "00100000",
                     238 => "10010111",
                     239 => "10001111",
                     240 => "10101101",
                     241 => "01110110",
                     242 => "00000111",
                     243 => "01001010",
                     244 => "10110000",
                     245 => "00100101",
                     246 => "10101101",
                     247 => "01000111",
                     248 => "00000111",
                     249 => "11110000",
                     250 => "00000101",
                     251 => "11001110",
                     252 => "01000111",
                     253 => "00000111",
                     254 => "11010000",
                     255 => "00011001",
                     256 => "10100010",
                     257 => "00010100",
                     258 => "11001110",
                     259 => "01111111",
                     260 => "00000111",
                     261 => "00010000",
                     262 => "00000111",
                     263 => "10101001",
                     264 => "00010001",
                     265 => "10001101",
                     266 => "01111111",
                     267 => "00000111",
                     268 => "10100010",
                     269 => "00100011",
                     270 => "10111101",
                     271 => "10000000",
                     272 => "00000111",
                     273 => "11110000",
                     274 => "00000011",
                     275 => "11011110",
                     276 => "10000000",
                     277 => "00000111",
                     278 => "11001010",
                     279 => "00010000",
                     280 => "11110101",
                     281 => "11100110",
                     282 => "00001001",
                     283 => "10100010",
                     284 => "00000000",
                     285 => "10100000",
                     286 => "00000111",
                     287 => "10101101",
                     288 => "10100111",
                     289 => "00000111",
                     290 => "00101001",
                     291 => "00000010",
                     292 => "10000101",
                     293 => "00000000",
                     294 => "10101101",
                     295 => "10101000",
                     296 => "00000111",
                     297 => "00101001",
                     298 => "00000010",
                     299 => "01000101",
                     300 => "00000000",
                     301 => "00011000",
                     302 => "11110000",
                     303 => "00000001",
                     304 => "00111000",
                     305 => "01111110",
                     306 => "10100111",
                     307 => "00000111",
                     308 => "11101000",
                     309 => "10001000",
                     310 => "11010000",
                     311 => "11111001",
                     312 => "10101101",
                     313 => "00100010",
                     314 => "00000111",
                     315 => "11110000",
                     316 => "00011111",
                     317 => "10101101",
                     318 => "00000010",
                     319 => "00100000",
                     320 => "00101001",
                     321 => "01000000",
                     322 => "11010000",
                     323 => "11111001",
                     324 => "10101101",
                     325 => "01110110",
                     326 => "00000111",
                     327 => "01001010",
                     328 => "10110000",
                     329 => "00000110",
                     330 => "00100000",
                     331 => "00100011",
                     332 => "10000010",
                     333 => "00100000",
                     334 => "11000110",
                     335 => "10000001",
                     336 => "10101101",
                     337 => "00000010",
                     338 => "00100000",
                     339 => "00101001",
                     340 => "01000000",
                     341 => "11110000",
                     342 => "11111001",
                     343 => "10100000",
                     344 => "00010100",
                     345 => "10001000",
                     346 => "11010000",
                     347 => "11111101",
                     348 => "10101101",
                     349 => "00111111",
                     350 => "00000111",
                     351 => "10001101",
                     352 => "00000101",
                     353 => "00100000",
                     354 => "10101101",
                     355 => "01000000",
                     356 => "00000111",
                     357 => "10001101",
                     358 => "00000101",
                     359 => "00100000",
                     360 => "10101101",
                     361 => "01111000",
                     362 => "00000111",
                     363 => "01001000",
                     364 => "10001101",
                     365 => "00000000",
                     366 => "00100000",
                     367 => "10101101",
                     368 => "01110110",
                     369 => "00000111",
                     370 => "01001010",
                     371 => "10110000",
                     372 => "00000011",
                     373 => "00100000",
                     374 => "00010010",
                     375 => "10000010",
                     376 => "10101101",
                     377 => "00000010",
                     378 => "00100000",
                     379 => "01101000",
                     380 => "00001001",
                     381 => "10000000",
                     382 => "10001101",
                     383 => "00000000",
                     384 => "00100000",
                     385 => "01000000",
                     386 => "10101101",
                     387 => "01110000",
                     388 => "00000111",
                     389 => "11001001",
                     390 => "00000010",
                     391 => "11110000",
                     392 => "00001011",
                     393 => "11001001",
                     394 => "00000001",
                     395 => "11010000",
                     396 => "00111000",
                     397 => "10101101",
                     398 => "01110010",
                     399 => "00000111",
                     400 => "11001001",
                     401 => "00000011",
                     402 => "11010000",
                     403 => "00110001",
                     404 => "10101101",
                     405 => "01110111",
                     406 => "00000111",
                     407 => "11110000",
                     408 => "00000100",
                     409 => "11001110",
                     410 => "01110111",
                     411 => "00000111",
                     412 => "01100000",
                     413 => "10101101",
                     414 => "11111100",
                     415 => "00000110",
                     416 => "00101001",
                     417 => "00010000",
                     418 => "11110000",
                     419 => "00011001",
                     420 => "10101101",
                     421 => "01110110",
                     422 => "00000111",
                     423 => "00101001",
                     424 => "10000000",
                     425 => "11010000",
                     426 => "00011010",
                     427 => "10101001",
                     428 => "00101011",
                     429 => "10001101",
                     430 => "01110111",
                     431 => "00000111",
                     432 => "10101101",
                     433 => "01110110",
                     434 => "00000111",
                     435 => "10101000",
                     436 => "11001000",
                     437 => "10000100",
                     438 => "11111010",
                     439 => "01001001",
                     440 => "00000001",
                     441 => "00001001",
                     442 => "10000000",
                     443 => "11010000",
                     444 => "00000101",
                     445 => "10101101",
                     446 => "01110110",
                     447 => "00000111",
                     448 => "00101001",
                     449 => "01111111",
                     450 => "10001101",
                     451 => "01110110",
                     452 => "00000111",
                     453 => "01100000",
                     454 => "10101100",
                     455 => "01001110",
                     456 => "00000111",
                     457 => "10101001",
                     458 => "00101000",
                     459 => "10000101",
                     460 => "00000000",
                     461 => "10100010",
                     462 => "00001110",
                     463 => "10111101",
                     464 => "11100100",
                     465 => "00000110",
                     466 => "11000101",
                     467 => "00000000",
                     468 => "10010000",
                     469 => "00001111",
                     470 => "10101100",
                     471 => "11100000",
                     472 => "00000110",
                     473 => "00011000",
                     474 => "01111001",
                     475 => "11100001",
                     476 => "00000110",
                     477 => "10010000",
                     478 => "00000011",
                     479 => "00011000",
                     480 => "01100101",
                     481 => "00000000",
                     482 => "10011101",
                     483 => "11100100",
                     484 => "00000110",
                     485 => "11001010",
                     486 => "00010000",
                     487 => "11100111",
                     488 => "10101110",
                     489 => "11100000",
                     490 => "00000110",
                     491 => "11101000",
                     492 => "11100000",
                     493 => "00000011",
                     494 => "11010000",
                     495 => "00000010",
                     496 => "10100010",
                     497 => "00000000",
                     498 => "10001110",
                     499 => "11100000",
                     500 => "00000110",
                     501 => "10100010",
                     502 => "00001000",
                     503 => "10100000",
                     504 => "00000010",
                     505 => "10111001",
                     506 => "11101001",
                     507 => "00000110",
                     508 => "10011101",
                     509 => "11110001",
                     510 => "00000110",
                     511 => "00011000",
                     512 => "01101001",
                     513 => "00001000",
                     514 => "10011101",
                     515 => "11110010",
                     516 => "00000110",
                     517 => "00011000",
                     518 => "01101001",
                     519 => "00001000",
                     520 => "10011101",
                     521 => "11110011",
                     522 => "00000110",
                     523 => "11001010",
                     524 => "11001010",
                     525 => "11001010",
                     526 => "10001000",
                     527 => "00010000",
                     528 => "11101000",
                     529 => "01100000",
                     530 => "10101101",
                     531 => "01110000",
                     532 => "00000111",
                     533 => "00100000",
                     534 => "00000100",
                     535 => "10001110",
                     536 => "00110001",
                     537 => "10000010",
                     538 => "11011100",
                     539 => "10101110",
                     540 => "10001011",
                     541 => "10000011",
                     542 => "00011000",
                     543 => "10010010",
                     544 => "10100000",
                     545 => "00000000",
                     546 => "00101100",
                     547 => "10100000",
                     548 => "00000100",
                     549 => "10101001",
                     550 => "11111000",
                     551 => "10011001",
                     552 => "00000000",
                     553 => "00000010",
                     554 => "11001000",
                     555 => "11001000",
                     556 => "11001000",
                     557 => "11001000",
                     558 => "11010000",
                     559 => "11110111",
                     560 => "01100000",
                     561 => "10101101",
                     562 => "01110010",
                     563 => "00000111",
                     564 => "00100000",
                     565 => "00000100",
                     566 => "10001110",
                     567 => "11001111",
                     568 => "10001111",
                     569 => "01100111",
                     570 => "10000101",
                     571 => "01100001",
                     572 => "10010000",
                     573 => "01000101",
                     574 => "10000010",
                     575 => "00000100",
                     576 => "00100000",
                     577 => "01110011",
                     578 => "00000001",
                     579 => "00000000",
                     580 => "00000000",
                     581 => "10100000",
                     582 => "00000000",
                     583 => "10101101",
                     584 => "11111100",
                     585 => "00000110",
                     586 => "00001101",
                     587 => "11111101",
                     588 => "00000110",
                     589 => "11001001",
                     590 => "00010000",
                     591 => "11110000",
                     592 => "00000100",
                     593 => "11001001",
                     594 => "10010000",
                     595 => "11010000",
                     596 => "00000011",
                     597 => "01001100",
                     598 => "11011000",
                     599 => "10000010",
                     600 => "11001001",
                     601 => "00100000",
                     602 => "11110000",
                     603 => "00011010",
                     604 => "10101110",
                     605 => "10100010",
                     606 => "00000111",
                     607 => "11010000",
                     608 => "00001011",
                     609 => "10001101",
                     610 => "10000000",
                     611 => "00000111",
                     612 => "00100000",
                     613 => "01101011",
                     614 => "10000011",
                     615 => "10110000",
                     616 => "01100000",
                     617 => "01001100",
                     618 => "11000000",
                     619 => "10000010",
                     620 => "10101110",
                     621 => "11111100",
                     622 => "00000111",
                     623 => "11110000",
                     624 => "01001010",
                     625 => "11001001",
                     626 => "01000000",
                     627 => "11010000",
                     628 => "01000110",
                     629 => "11001000",
                     630 => "10101101",
                     631 => "10100010",
                     632 => "00000111",
                     633 => "11110000",
                     634 => "01001110",
                     635 => "10101001",
                     636 => "00011000",
                     637 => "10001101",
                     638 => "10100010",
                     639 => "00000111",
                     640 => "10101101",
                     641 => "10000000",
                     642 => "00000111",
                     643 => "11010000",
                     644 => "00110110",
                     645 => "10101001",
                     646 => "00010000",
                     647 => "10001101",
                     648 => "10000000",
                     649 => "00000111",
                     650 => "11000000",
                     651 => "00000001",
                     652 => "11110000",
                     653 => "00001110",
                     654 => "10101101",
                     655 => "01111010",
                     656 => "00000111",
                     657 => "01001001",
                     658 => "00000001",
                     659 => "10001101",
                     660 => "01111010",
                     661 => "00000111",
                     662 => "00100000",
                     663 => "00100101",
                     664 => "10000011",
                     665 => "01001100",
                     666 => "10111011",
                     667 => "10000010",
                     668 => "10101110",
                     669 => "01101011",
                     670 => "00000111",
                     671 => "11101000",
                     672 => "10001010",
                     673 => "00101001",
                     674 => "00000111",
                     675 => "10001101",
                     676 => "01101011",
                     677 => "00000111",
                     678 => "00100000",
                     679 => "00001110",
                     680 => "10000011",
                     681 => "10111101",
                     682 => "00111111",
                     683 => "10000010",
                     684 => "10011101",
                     685 => "00000000",
                     686 => "00000011",
                     687 => "11101000",
                     688 => "11100000",
                     689 => "00000110",
                     690 => "00110000",
                     691 => "11110101",
                     692 => "10101100",
                     693 => "01011111",
                     694 => "00000111",
                     695 => "11001000",
                     696 => "10001100",
                     697 => "00000100",
                     698 => "00000011",
                     699 => "10101001",
                     700 => "00000000",
                     701 => "10001101",
                     702 => "11111100",
                     703 => "00000110",
                     704 => "00100000",
                     705 => "11101010",
                     706 => "10101110",
                     707 => "10100101",
                     708 => "00001110",
                     709 => "11001001",
                     710 => "00000110",
                     711 => "11010000",
                     712 => "01000100",
                     713 => "10101001",
                     714 => "00000000",
                     715 => "10001101",
                     716 => "01110000",
                     717 => "00000111",
                     718 => "10001101",
                     719 => "01110010",
                     720 => "00000111",
                     721 => "10001101",
                     722 => "00100010",
                     723 => "00000111",
                     724 => "11101110",
                     725 => "01110100",
                     726 => "00000111",
                     727 => "01100000",
                     728 => "10101100",
                     729 => "10100010",
                     730 => "00000111",
                     731 => "11110000",
                     732 => "11101100",
                     733 => "00001010",
                     734 => "10010000",
                     735 => "00000110",
                     736 => "10101101",
                     737 => "11111101",
                     738 => "00000111",
                     739 => "00100000",
                     740 => "00001110",
                     741 => "10000011",
                     742 => "00100000",
                     743 => "00000011",
                     744 => "10011100",
                     745 => "11101110",
                     746 => "01011101",
                     747 => "00000111",
                     748 => "11101110",
                     749 => "01100100",
                     750 => "00000111",
                     751 => "11101110",
                     752 => "01010111",
                     753 => "00000111",
                     754 => "11101110",
                     755 => "01110000",
                     756 => "00000111",
                     757 => "10101101",
                     758 => "11111100",
                     759 => "00000111",
                     760 => "10001101",
                     761 => "01101010",
                     762 => "00000111",
                     763 => "10101001",
                     764 => "00000000",
                     765 => "10001101",
                     766 => "01110010",
                     767 => "00000111",
                     768 => "10001101",
                     769 => "10100010",
                     770 => "00000111",
                     771 => "10100010",
                     772 => "00010111",
                     773 => "10101001",
                     774 => "00000000",
                     775 => "10011101",
                     776 => "11011101",
                     777 => "00000111",
                     778 => "11001010",
                     779 => "00010000",
                     780 => "11111010",
                     781 => "01100000",
                     782 => "10001101",
                     783 => "01011111",
                     784 => "00000111",
                     785 => "10001101",
                     786 => "01100110",
                     787 => "00000111",
                     788 => "10100010",
                     789 => "00000000",
                     790 => "10001110",
                     791 => "01100000",
                     792 => "00000111",
                     793 => "10001110",
                     794 => "01100111",
                     795 => "00000111",
                     796 => "01100000",
                     797 => "00000111",
                     798 => "00100010",
                     799 => "01001001",
                     800 => "10000011",
                     801 => "11001110",
                     802 => "00100100",
                     803 => "00100100",
                     804 => "00000000",
                     805 => "10100000",
                     806 => "00000111",
                     807 => "10111001",
                     808 => "00011101",
                     809 => "10000011",
                     810 => "10011001",
                     811 => "00000000",
                     812 => "00000011",
                     813 => "10001000",
                     814 => "00010000",
                     815 => "11110111",
                     816 => "10101101",
                     817 => "01111010",
                     818 => "00000111",
                     819 => "11110000",
                     820 => "00001010",
                     821 => "10101001",
                     822 => "00100100",
                     823 => "10001101",
                     824 => "00000100",
                     825 => "00000011",
                     826 => "10101001",
                     827 => "11001110",
                     828 => "10001101",
                     829 => "00000110",
                     830 => "00000011",
                     831 => "01100000",
                     832 => "00000001",
                     833 => "10000000",
                     834 => "00000010",
                     835 => "10000001",
                     836 => "01000001",
                     837 => "10000000",
                     838 => "00000001",
                     839 => "01000010",
                     840 => "11000010",
                     841 => "00000010",
                     842 => "10000000",
                     843 => "01000001",
                     844 => "11000001",
                     845 => "01000001",
                     846 => "11000001",
                     847 => "00000001",
                     848 => "11000001",
                     849 => "00000001",
                     850 => "00000010",
                     851 => "10000000",
                     852 => "00000000",
                     853 => "10011011",
                     854 => "00010000",
                     855 => "00011000",
                     856 => "00000101",
                     857 => "00101100",
                     858 => "00100000",
                     859 => "00100100",
                     860 => "00010101",
                     861 => "01011010",
                     862 => "00010000",
                     863 => "00100000",
                     864 => "00101000",
                     865 => "00110000",
                     866 => "00100000",
                     867 => "00010000",
                     868 => "10000000",
                     869 => "00100000",
                     870 => "00110000",
                     871 => "00110000",
                     872 => "00000001",
                     873 => "11111111",
                     874 => "00000000",
                     875 => "10101110",
                     876 => "00010111",
                     877 => "00000111",
                     878 => "10101101",
                     879 => "00011000",
                     880 => "00000111",
                     881 => "11010000",
                     882 => "00001101",
                     883 => "11101000",
                     884 => "11101110",
                     885 => "00010111",
                     886 => "00000111",
                     887 => "00111000",
                     888 => "10111101",
                     889 => "01010100",
                     890 => "10000011",
                     891 => "10001101",
                     892 => "00011000",
                     893 => "00000111",
                     894 => "11110000",
                     895 => "00001010",
                     896 => "10111101",
                     897 => "00111111",
                     898 => "10000011",
                     899 => "10001101",
                     900 => "11111100",
                     901 => "00000110",
                     902 => "11001110",
                     903 => "00011000",
                     904 => "00000111",
                     905 => "00011000",
                     906 => "01100000",
                     907 => "00100000",
                     908 => "10100000",
                     909 => "10000011",
                     910 => "10101101",
                     911 => "01110010",
                     912 => "00000111",
                     913 => "11110000",
                     914 => "00000111",
                     915 => "10100010",
                     916 => "00000000",
                     917 => "10000110",
                     918 => "00001000",
                     919 => "00100000",
                     920 => "01001101",
                     921 => "11000000",
                     922 => "00100000",
                     923 => "00110001",
                     924 => "11110001",
                     925 => "01001100",
                     926 => "11110000",
                     927 => "11101110",
                     928 => "10101101",
                     929 => "01110010",
                     930 => "00000111",
                     931 => "00100000",
                     932 => "00000100",
                     933 => "10001110",
                     934 => "10110100",
                     935 => "11001111",
                     936 => "10110000",
                     937 => "10000011",
                     938 => "10111101",
                     939 => "10000011",
                     940 => "11110110",
                     941 => "10000011",
                     942 => "01100001",
                     943 => "10000100",
                     944 => "10101110",
                     945 => "00011011",
                     946 => "00000111",
                     947 => "11101000",
                     948 => "10000110",
                     949 => "00110100",
                     950 => "10101001",
                     951 => "00001000",
                     952 => "10000101",
                     953 => "11111100",
                     954 => "01001100",
                     955 => "01001110",
                     956 => "10000111",
                     957 => "10100000",
                     958 => "00000000",
                     959 => "10000100",
                     960 => "00110101",
                     961 => "10100101",
                     962 => "01101101",
                     963 => "11000101",
                     964 => "00110100",
                     965 => "11010000",
                     966 => "00000110",
                     967 => "10100101",
                     968 => "10000110",
                     969 => "11001001",
                     970 => "01100000",
                     971 => "10110000",
                     972 => "00000011",
                     973 => "11100110",
                     974 => "00110101",
                     975 => "11001000",
                     976 => "10011000",
                     977 => "00100000",
                     978 => "11100110",
                     979 => "10110000",
                     980 => "10101101",
                     981 => "00011010",
                     982 => "00000111",
                     983 => "11000101",
                     984 => "00110100",
                     985 => "11110000",
                     986 => "00010110",
                     987 => "10101101",
                     988 => "01101000",
                     989 => "00000111",
                     990 => "00011000",
                     991 => "01101001",
                     992 => "10000000",
                     993 => "10001101",
                     994 => "01101000",
                     995 => "00000111",
                     996 => "10101001",
                     997 => "00000001",
                     998 => "01101001",
                     999 => "00000000",
                     1000 => "10101000",
                     1001 => "00100000",
                     1002 => "11000100",
                     1003 => "10101111",
                     1004 => "00100000",
                     1005 => "01101111",
                     1006 => "10101111",
                     1007 => "11100110",
                     1008 => "00110101",
                     1009 => "10100101",
                     1010 => "00110101",
                     1011 => "11110000",
                     1012 => "01101000",
                     1013 => "01100000",
                     1014 => "10101101",
                     1015 => "01001001",
                     1016 => "00000111",
                     1017 => "11010000",
                     1018 => "01001000",
                     1019 => "10101101",
                     1020 => "00011001",
                     1021 => "00000111",
                     1022 => "11110000",
                     1023 => "00011000",
                     1024 => "11001001",
                     1025 => "00001001",
                     1026 => "10110000",
                     1027 => "00111111",
                     1028 => "10101100",
                     1029 => "01011111",
                     1030 => "00000111",
                     1031 => "11000000",
                     1032 => "00000111",
                     1033 => "11010000",
                     1034 => "00001001",
                     1035 => "11001001",
                     1036 => "00000011",
                     1037 => "10010000",
                     1038 => "00110100",
                     1039 => "11101001",
                     1040 => "00000001",
                     1041 => "01001100",
                     1042 => "00011000",
                     1043 => "10000100",
                     1044 => "11001001",
                     1045 => "00000010",
                     1046 => "10010000",
                     1047 => "00101011",
                     1048 => "10101000",
                     1049 => "11010000",
                     1050 => "00001000",
                     1051 => "10101101",
                     1052 => "01010011",
                     1053 => "00000111",
                     1054 => "11110000",
                     1055 => "00010100",
                     1056 => "11001000",
                     1057 => "11010000",
                     1058 => "00010001",
                     1059 => "11001000",
                     1060 => "10101101",
                     1061 => "01011111",
                     1062 => "00000111",
                     1063 => "11001001",
                     1064 => "00000111",
                     1065 => "11110000",
                     1066 => "00001001",
                     1067 => "10001000",
                     1068 => "11000000",
                     1069 => "00000100",
                     1070 => "10110000",
                     1071 => "00100110",
                     1072 => "11000000",
                     1073 => "00000011",
                     1074 => "10110000",
                     1075 => "00001111",
                     1076 => "11000000",
                     1077 => "00000011",
                     1078 => "11010000",
                     1079 => "00000100",
                     1080 => "10101001",
                     1081 => "00000100",
                     1082 => "10000101",
                     1083 => "11111100",
                     1084 => "10011000",
                     1085 => "00011000",
                     1086 => "01101001",
                     1087 => "00001100",
                     1088 => "10001101",
                     1089 => "01110011",
                     1090 => "00000111",
                     1091 => "10101101",
                     1092 => "01001001",
                     1093 => "00000111",
                     1094 => "00011000",
                     1095 => "01101001",
                     1096 => "00000100",
                     1097 => "10001101",
                     1098 => "01001001",
                     1099 => "00000111",
                     1100 => "10101101",
                     1101 => "00011001",
                     1102 => "00000111",
                     1103 => "01101001",
                     1104 => "00000000",
                     1105 => "10001101",
                     1106 => "00011001",
                     1107 => "00000111",
                     1108 => "11001001",
                     1109 => "00000111",
                     1110 => "10010000",
                     1111 => "00001000",
                     1112 => "10101001",
                     1113 => "00000110",
                     1114 => "10001101",
                     1115 => "10100001",
                     1116 => "00000111",
                     1117 => "11101110",
                     1118 => "01110010",
                     1119 => "00000111",
                     1120 => "01100000",
                     1121 => "10101101",
                     1122 => "10100001",
                     1123 => "00000111",
                     1124 => "11010000",
                     1125 => "00100000",
                     1126 => "10101100",
                     1127 => "01011111",
                     1128 => "00000111",
                     1129 => "11000000",
                     1130 => "00000111",
                     1131 => "10110000",
                     1132 => "00011010",
                     1133 => "10101001",
                     1134 => "00000000",
                     1135 => "10001101",
                     1136 => "01100000",
                     1137 => "00000111",
                     1138 => "10001101",
                     1139 => "01011100",
                     1140 => "00000111",
                     1141 => "10001101",
                     1142 => "01110010",
                     1143 => "00000111",
                     1144 => "11101110",
                     1145 => "01011111",
                     1146 => "00000111",
                     1147 => "00100000",
                     1148 => "00000011",
                     1149 => "10011100",
                     1150 => "11101110",
                     1151 => "01010111",
                     1152 => "00000111",
                     1153 => "10101001",
                     1154 => "00000001",
                     1155 => "10001101",
                     1156 => "01110000",
                     1157 => "00000111",
                     1158 => "01100000",
                     1159 => "10101101",
                     1160 => "11111100",
                     1161 => "00000110",
                     1162 => "00001101",
                     1163 => "11111101",
                     1164 => "00000110",
                     1165 => "00101001",
                     1166 => "01000000",
                     1167 => "11110000",
                     1168 => "00001101",
                     1169 => "10101001",
                     1170 => "00000001",
                     1171 => "10001101",
                     1172 => "11111100",
                     1173 => "00000111",
                     1174 => "10101001",
                     1175 => "11111111",
                     1176 => "10001101",
                     1177 => "01011010",
                     1178 => "00000111",
                     1179 => "00100000",
                     1180 => "01001000",
                     1181 => "10010010",
                     1182 => "01100000",
                     1183 => "11111111",
                     1184 => "11111111",
                     1185 => "11110110",
                     1186 => "11111011",
                     1187 => "11110111",
                     1188 => "11111011",
                     1189 => "11111000",
                     1190 => "11111011",
                     1191 => "11111001",
                     1192 => "11111011",
                     1193 => "11111010",
                     1194 => "11111011",
                     1195 => "11110110",
                     1196 => "01010000",
                     1197 => "11110111",
                     1198 => "01010000",
                     1199 => "11111000",
                     1200 => "01010000",
                     1201 => "11111001",
                     1202 => "01010000",
                     1203 => "11111010",
                     1204 => "01010000",
                     1205 => "11111101",
                     1206 => "11111110",
                     1207 => "11111111",
                     1208 => "01000001",
                     1209 => "01000010",
                     1210 => "01000100",
                     1211 => "01000101",
                     1212 => "01001000",
                     1213 => "00110001",
                     1214 => "00110010",
                     1215 => "00110100",
                     1216 => "00110101",
                     1217 => "00111000",
                     1218 => "00000000",
                     1219 => "10111101",
                     1220 => "00010000",
                     1221 => "00000001",
                     1222 => "11110000",
                     1223 => "10111110",
                     1224 => "11001001",
                     1225 => "00001011",
                     1226 => "10010000",
                     1227 => "00000101",
                     1228 => "10101001",
                     1229 => "00001011",
                     1230 => "10011101",
                     1231 => "00010000",
                     1232 => "00000001",
                     1233 => "10101000",
                     1234 => "10111101",
                     1235 => "00101100",
                     1236 => "00000001",
                     1237 => "11010000",
                     1238 => "00000100",
                     1239 => "10011101",
                     1240 => "00010000",
                     1241 => "00000001",
                     1242 => "01100000",
                     1243 => "11011110",
                     1244 => "00101100",
                     1245 => "00000001",
                     1246 => "11001001",
                     1247 => "00101011",
                     1248 => "11010000",
                     1249 => "00011110",
                     1250 => "11000000",
                     1251 => "00001011",
                     1252 => "11010000",
                     1253 => "00000111",
                     1254 => "11101110",
                     1255 => "01011010",
                     1256 => "00000111",
                     1257 => "10101001",
                     1258 => "01000000",
                     1259 => "10000101",
                     1260 => "11111110",
                     1261 => "10111001",
                     1262 => "10110111",
                     1263 => "10000100",
                     1264 => "01001010",
                     1265 => "01001010",
                     1266 => "01001010",
                     1267 => "01001010",
                     1268 => "10101010",
                     1269 => "10111001",
                     1270 => "10110111",
                     1271 => "10000100",
                     1272 => "00101001",
                     1273 => "00001111",
                     1274 => "10011101",
                     1275 => "00110100",
                     1276 => "00000001",
                     1277 => "00100000",
                     1278 => "00101100",
                     1279 => "10111100",
                     1280 => "10111100",
                     1281 => "11100101",
                     1282 => "00000110",
                     1283 => "10110101",
                     1284 => "00010110",
                     1285 => "11001001",
                     1286 => "00010010",
                     1287 => "11110000",
                     1288 => "00100010",
                     1289 => "11001001",
                     1290 => "00001101",
                     1291 => "11110000",
                     1292 => "00011110",
                     1293 => "11001001",
                     1294 => "00000101",
                     1295 => "11110000",
                     1296 => "00010010",
                     1297 => "11001001",
                     1298 => "00001010",
                     1299 => "11110000",
                     1300 => "00010110",
                     1301 => "11001001",
                     1302 => "00001011",
                     1303 => "11110000",
                     1304 => "00010010",
                     1305 => "11001001",
                     1306 => "00001001",
                     1307 => "10110000",
                     1308 => "00000110",
                     1309 => "10110101",
                     1310 => "00011110",
                     1311 => "11001001",
                     1312 => "00000010",
                     1313 => "10110000",
                     1314 => "00001000",
                     1315 => "10101110",
                     1316 => "11101110",
                     1317 => "00000011",
                     1318 => "10111100",
                     1319 => "11101100",
                     1320 => "00000110",
                     1321 => "10100110",
                     1322 => "00001000",
                     1323 => "10111101",
                     1324 => "00011110",
                     1325 => "00000001",
                     1326 => "11001001",
                     1327 => "00011000",
                     1328 => "10010000",
                     1329 => "00000101",
                     1330 => "11101001",
                     1331 => "00000001",
                     1332 => "10011101",
                     1333 => "00011110",
                     1334 => "00000001",
                     1335 => "10111101",
                     1336 => "00011110",
                     1337 => "00000001",
                     1338 => "11101001",
                     1339 => "00001000",
                     1340 => "00100000",
                     1341 => "11001000",
                     1342 => "11100101",
                     1343 => "10111101",
                     1344 => "00010111",
                     1345 => "00000001",
                     1346 => "10011001",
                     1347 => "00000011",
                     1348 => "00000010",
                     1349 => "00011000",
                     1350 => "01101001",
                     1351 => "00001000",
                     1352 => "10011001",
                     1353 => "00000111",
                     1354 => "00000010",
                     1355 => "10101001",
                     1356 => "00000010",
                     1357 => "10011001",
                     1358 => "00000010",
                     1359 => "00000010",
                     1360 => "10011001",
                     1361 => "00000110",
                     1362 => "00000010",
                     1363 => "10111101",
                     1364 => "00010000",
                     1365 => "00000001",
                     1366 => "00001010",
                     1367 => "10101010",
                     1368 => "10111101",
                     1369 => "10011111",
                     1370 => "10000100",
                     1371 => "10011001",
                     1372 => "00000001",
                     1373 => "00000010",
                     1374 => "10111101",
                     1375 => "10100000",
                     1376 => "10000100",
                     1377 => "10011001",
                     1378 => "00000101",
                     1379 => "00000010",
                     1380 => "10100110",
                     1381 => "00001000",
                     1382 => "01100000",
                     1383 => "10101101",
                     1384 => "00111100",
                     1385 => "00000111",
                     1386 => "00100000",
                     1387 => "00000100",
                     1388 => "10001110",
                     1389 => "10001011",
                     1390 => "10000101",
                     1391 => "10011011",
                     1392 => "10000101",
                     1393 => "01010010",
                     1394 => "10000110",
                     1395 => "01011010",
                     1396 => "10000110",
                     1397 => "10010011",
                     1398 => "10000110",
                     1399 => "10011101",
                     1400 => "10001000",
                     1401 => "10101000",
                     1402 => "10000110",
                     1403 => "10011101",
                     1404 => "10001000",
                     1405 => "11100110",
                     1406 => "10000110",
                     1407 => "10111111",
                     1408 => "10000101",
                     1409 => "11100011",
                     1410 => "10000101",
                     1411 => "01000011",
                     1412 => "10000110",
                     1413 => "11111111",
                     1414 => "10000110",
                     1415 => "00110010",
                     1416 => "10000111",
                     1417 => "01001001",
                     1418 => "10000111",
                     1419 => "00100000",
                     1420 => "00100000",
                     1421 => "10000010",
                     1422 => "00100000",
                     1423 => "00011001",
                     1424 => "10001110",
                     1425 => "10101101",
                     1426 => "01110000",
                     1427 => "00000111",
                     1428 => "11110000",
                     1429 => "00110010",
                     1430 => "10100010",
                     1431 => "00000011",
                     1432 => "01001100",
                     1433 => "11000101",
                     1434 => "10000101",
                     1435 => "10101101",
                     1436 => "01000100",
                     1437 => "00000111",
                     1438 => "01001000",
                     1439 => "10101101",
                     1440 => "01010110",
                     1441 => "00000111",
                     1442 => "01001000",
                     1443 => "10101001",
                     1444 => "00000000",
                     1445 => "10001101",
                     1446 => "01010110",
                     1447 => "00000111",
                     1448 => "10101001",
                     1449 => "00000010",
                     1450 => "10001101",
                     1451 => "01000100",
                     1452 => "00000111",
                     1453 => "00100000",
                     1454 => "11110001",
                     1455 => "10000101",
                     1456 => "01101000",
                     1457 => "10001101",
                     1458 => "01010110",
                     1459 => "00000111",
                     1460 => "01101000",
                     1461 => "10001101",
                     1462 => "01000100",
                     1463 => "00000111",
                     1464 => "01001100",
                     1465 => "01000101",
                     1466 => "10000111",
                     1467 => "00000001",
                     1468 => "00000010",
                     1469 => "00000011",
                     1470 => "00000100",
                     1471 => "10101100",
                     1472 => "01001110",
                     1473 => "00000111",
                     1474 => "10111110",
                     1475 => "10111011",
                     1476 => "10000101",
                     1477 => "10001110",
                     1478 => "01110011",
                     1479 => "00000111",
                     1480 => "01001100",
                     1481 => "01000101",
                     1482 => "10000111",
                     1483 => "00000000",
                     1484 => "00001001",
                     1485 => "00001010",
                     1486 => "00000100",
                     1487 => "00100010",
                     1488 => "00100010",
                     1489 => "00001111",
                     1490 => "00001111",
                     1491 => "00001111",
                     1492 => "00100010",
                     1493 => "00001111",
                     1494 => "00001111",
                     1495 => "00100010",
                     1496 => "00010110",
                     1497 => "00100111",
                     1498 => "00011000",
                     1499 => "00100010",
                     1500 => "00110000",
                     1501 => "00100111",
                     1502 => "00011001",
                     1503 => "00100010",
                     1504 => "00110111",
                     1505 => "00100111",
                     1506 => "00010110",
                     1507 => "10101100",
                     1508 => "01000100",
                     1509 => "00000111",
                     1510 => "11110000",
                     1511 => "00000110",
                     1512 => "10111001",
                     1513 => "11000111",
                     1514 => "10000101",
                     1515 => "10001101",
                     1516 => "01110011",
                     1517 => "00000111",
                     1518 => "11101110",
                     1519 => "00111100",
                     1520 => "00000111",
                     1521 => "10101110",
                     1522 => "00000000",
                     1523 => "00000011",
                     1524 => "10100000",
                     1525 => "00000000",
                     1526 => "10101101",
                     1527 => "01010011",
                     1528 => "00000111",
                     1529 => "11110000",
                     1530 => "00000010",
                     1531 => "10100000",
                     1532 => "00000100",
                     1533 => "10101101",
                     1534 => "01010110",
                     1535 => "00000111",
                     1536 => "11001001",
                     1537 => "00000010",
                     1538 => "11010000",
                     1539 => "00000010",
                     1540 => "10100000",
                     1541 => "00001000",
                     1542 => "10101001",
                     1543 => "00000011",
                     1544 => "10000101",
                     1545 => "00000000",
                     1546 => "10111001",
                     1547 => "11010111",
                     1548 => "10000101",
                     1549 => "10011101",
                     1550 => "00000100",
                     1551 => "00000011",
                     1552 => "11001000",
                     1553 => "11101000",
                     1554 => "11000110",
                     1555 => "00000000",
                     1556 => "00010000",
                     1557 => "11110100",
                     1558 => "10101110",
                     1559 => "00000000",
                     1560 => "00000011",
                     1561 => "10101100",
                     1562 => "01000100",
                     1563 => "00000111",
                     1564 => "11010000",
                     1565 => "00000011",
                     1566 => "10101100",
                     1567 => "01001110",
                     1568 => "00000111",
                     1569 => "10111001",
                     1570 => "11001111",
                     1571 => "10000101",
                     1572 => "10011101",
                     1573 => "00000100",
                     1574 => "00000011",
                     1575 => "10101001",
                     1576 => "00111111",
                     1577 => "10011101",
                     1578 => "00000001",
                     1579 => "00000011",
                     1580 => "10101001",
                     1581 => "00010000",
                     1582 => "10011101",
                     1583 => "00000010",
                     1584 => "00000011",
                     1585 => "10101001",
                     1586 => "00000100",
                     1587 => "10011101",
                     1588 => "00000011",
                     1589 => "00000011",
                     1590 => "10101001",
                     1591 => "00000000",
                     1592 => "10011101",
                     1593 => "00001000",
                     1594 => "00000011",
                     1595 => "10001010",
                     1596 => "00011000",
                     1597 => "01101001",
                     1598 => "00000111",
                     1599 => "10001101",
                     1600 => "00000000",
                     1601 => "00000011",
                     1602 => "01100000",
                     1603 => "10101101",
                     1604 => "00110011",
                     1605 => "00000111",
                     1606 => "11001001",
                     1607 => "00000001",
                     1608 => "11010000",
                     1609 => "00000101",
                     1610 => "10101001",
                     1611 => "00001011",
                     1612 => "10001101",
                     1613 => "01110011",
                     1614 => "00000111",
                     1615 => "01001100",
                     1616 => "01000101",
                     1617 => "10000111",
                     1618 => "10101001",
                     1619 => "00000000",
                     1620 => "00100000",
                     1621 => "00001000",
                     1622 => "10001000",
                     1623 => "01001100",
                     1624 => "01000101",
                     1625 => "10000111",
                     1626 => "00100000",
                     1627 => "00110101",
                     1628 => "10111100",
                     1629 => "10101110",
                     1630 => "00000000",
                     1631 => "00000011",
                     1632 => "10101001",
                     1633 => "00100000",
                     1634 => "10011101",
                     1635 => "00000001",
                     1636 => "00000011",
                     1637 => "10101001",
                     1638 => "01110011",
                     1639 => "10011101",
                     1640 => "00000010",
                     1641 => "00000011",
                     1642 => "10101001",
                     1643 => "00000011",
                     1644 => "10011101",
                     1645 => "00000011",
                     1646 => "00000011",
                     1647 => "10101100",
                     1648 => "01011111",
                     1649 => "00000111",
                     1650 => "11001000",
                     1651 => "10011000",
                     1652 => "10011101",
                     1653 => "00000100",
                     1654 => "00000011",
                     1655 => "10101001",
                     1656 => "00101000",
                     1657 => "10011101",
                     1658 => "00000101",
                     1659 => "00000011",
                     1660 => "10101100",
                     1661 => "01011100",
                     1662 => "00000111",
                     1663 => "11001000",
                     1664 => "10011000",
                     1665 => "10011101",
                     1666 => "00000110",
                     1667 => "00000011",
                     1668 => "10101001",
                     1669 => "00000000",
                     1670 => "10011101",
                     1671 => "00000111",
                     1672 => "00000011",
                     1673 => "10001010",
                     1674 => "00011000",
                     1675 => "01101001",
                     1676 => "00000110",
                     1677 => "10001101",
                     1678 => "00000000",
                     1679 => "00000011",
                     1680 => "01001100",
                     1681 => "01000101",
                     1682 => "10000111",
                     1683 => "10101101",
                     1684 => "01011001",
                     1685 => "00000111",
                     1686 => "11110000",
                     1687 => "00001010",
                     1688 => "10101001",
                     1689 => "00000000",
                     1690 => "10001101",
                     1691 => "01011001",
                     1692 => "00000111",
                     1693 => "10101001",
                     1694 => "00000010",
                     1695 => "01001100",
                     1696 => "11000111",
                     1697 => "10000110",
                     1698 => "11101110",
                     1699 => "00111100",
                     1700 => "00000111",
                     1701 => "01001100",
                     1702 => "01000101",
                     1703 => "10000111",
                     1704 => "10101101",
                     1705 => "01110000",
                     1706 => "00000111",
                     1707 => "11110000",
                     1708 => "00110011",
                     1709 => "11001001",
                     1710 => "00000011",
                     1711 => "11110000",
                     1712 => "00100010",
                     1713 => "10101101",
                     1714 => "01010010",
                     1715 => "00000111",
                     1716 => "11010000",
                     1717 => "00101010",
                     1718 => "10101100",
                     1719 => "01001110",
                     1720 => "00000111",
                     1721 => "11000000",
                     1722 => "00000011",
                     1723 => "11110000",
                     1724 => "00000101",
                     1725 => "10101101",
                     1726 => "01101001",
                     1727 => "00000111",
                     1728 => "11010000",
                     1729 => "00011110",
                     1730 => "00100000",
                     1731 => "10101011",
                     1732 => "11101111",
                     1733 => "10101001",
                     1734 => "00000001",
                     1735 => "00100000",
                     1736 => "00001000",
                     1737 => "10001000",
                     1738 => "00100000",
                     1739 => "10100101",
                     1740 => "10001000",
                     1741 => "10101001",
                     1742 => "00000000",
                     1743 => "10001101",
                     1744 => "01110100",
                     1745 => "00000111",
                     1746 => "01100000",
                     1747 => "10101001",
                     1748 => "00010010",
                     1749 => "10001101",
                     1750 => "10100000",
                     1751 => "00000111",
                     1752 => "10101001",
                     1753 => "00000011",
                     1754 => "00100000",
                     1755 => "00001000",
                     1756 => "10001000",
                     1757 => "01001100",
                     1758 => "01001110",
                     1759 => "10000111",
                     1760 => "10101001",
                     1761 => "00001000",
                     1762 => "10001101",
                     1763 => "00111100",
                     1764 => "00000111",
                     1765 => "01100000",
                     1766 => "11101110",
                     1767 => "01110100",
                     1768 => "00000111",
                     1769 => "00100000",
                     1770 => "10110000",
                     1771 => "10010010",
                     1772 => "10101101",
                     1773 => "00011111",
                     1774 => "00000111",
                     1775 => "11010000",
                     1776 => "11111000",
                     1777 => "11001110",
                     1778 => "00011110",
                     1779 => "00000111",
                     1780 => "00010000",
                     1781 => "00000011",
                     1782 => "11101110",
                     1783 => "00111100",
                     1784 => "00000111",
                     1785 => "10101001",
                     1786 => "00000110",
                     1787 => "10001101",
                     1788 => "01110011",
                     1789 => "00000111",
                     1790 => "01100000",
                     1791 => "10101101",
                     1792 => "01110000",
                     1793 => "00000111",
                     1794 => "11010000",
                     1795 => "01001010",
                     1796 => "10101001",
                     1797 => "00011110",
                     1798 => "10001101",
                     1799 => "00000110",
                     1800 => "00100000",
                     1801 => "10101001",
                     1802 => "11000000",
                     1803 => "10001101",
                     1804 => "00000110",
                     1805 => "00100000",
                     1806 => "10101001",
                     1807 => "00000011",
                     1808 => "10000101",
                     1809 => "00000001",
                     1810 => "10100000",
                     1811 => "00000000",
                     1812 => "10000100",
                     1813 => "00000000",
                     1814 => "10101101",
                     1815 => "00000111",
                     1816 => "00100000",
                     1817 => "10101101",
                     1818 => "00000111",
                     1819 => "00100000",
                     1820 => "10010001",
                     1821 => "00000000",
                     1822 => "11001000",
                     1823 => "11010000",
                     1824 => "00000010",
                     1825 => "11100110",
                     1826 => "00000001",
                     1827 => "10100101",
                     1828 => "00000001",
                     1829 => "11001001",
                     1830 => "00000100",
                     1831 => "11010000",
                     1832 => "11110000",
                     1833 => "11000000",
                     1834 => "00111010",
                     1835 => "10010000",
                     1836 => "11101100",
                     1837 => "10101001",
                     1838 => "00000101",
                     1839 => "01001100",
                     1840 => "01001100",
                     1841 => "10000110",
                     1842 => "10101101",
                     1843 => "01110000",
                     1844 => "00000111",
                     1845 => "11010000",
                     1846 => "00010111",
                     1847 => "10100010",
                     1848 => "00000000",
                     1849 => "10011101",
                     1850 => "00000000",
                     1851 => "00000011",
                     1852 => "10011101",
                     1853 => "00000000",
                     1854 => "00000100",
                     1855 => "11001010",
                     1856 => "11010000",
                     1857 => "11110111",
                     1858 => "00100000",
                     1859 => "00100101",
                     1860 => "10000011",
                     1861 => "11101110",
                     1862 => "00111100",
                     1863 => "00000111",
                     1864 => "01100000",
                     1865 => "10101001",
                     1866 => "11111010",
                     1867 => "00100000",
                     1868 => "00111011",
                     1869 => "10111100",
                     1870 => "11101110",
                     1871 => "01110010",
                     1872 => "00000111",
                     1873 => "01100000",
                     1874 => "00100000",
                     1875 => "01000011",
                     1876 => "00000101",
                     1877 => "00010110",
                     1878 => "00001010",
                     1879 => "00011011",
                     1880 => "00010010",
                     1881 => "00011000",
                     1882 => "00100000",
                     1883 => "01010010",
                     1884 => "00001011",
                     1885 => "00100000",
                     1886 => "00011000",
                     1887 => "00011011",
                     1888 => "00010101",
                     1889 => "00001101",
                     1890 => "00100100",
                     1891 => "00100100",
                     1892 => "00011101",
                     1893 => "00010010",
                     1894 => "00010110",
                     1895 => "00001110",
                     1896 => "00100000",
                     1897 => "01101000",
                     1898 => "00000101",
                     1899 => "00000000",
                     1900 => "00100100",
                     1901 => "00100100",
                     1902 => "00101110",
                     1903 => "00101001",
                     1904 => "00100011",
                     1905 => "11000000",
                     1906 => "01111111",
                     1907 => "10101010",
                     1908 => "00100011",
                     1909 => "11000010",
                     1910 => "00000001",
                     1911 => "11101010",
                     1912 => "11111111",
                     1913 => "00100001",
                     1914 => "11001101",
                     1915 => "00000111",
                     1916 => "00100100",
                     1917 => "00100100",
                     1918 => "00101001",
                     1919 => "00100100",
                     1920 => "00100100",
                     1921 => "00100100",
                     1922 => "00100100",
                     1923 => "00100001",
                     1924 => "01001011",
                     1925 => "00001001",
                     1926 => "00100000",
                     1927 => "00011000",
                     1928 => "00011011",
                     1929 => "00010101",
                     1930 => "00001101",
                     1931 => "00100100",
                     1932 => "00100100",
                     1933 => "00101000",
                     1934 => "00100100",
                     1935 => "00100010",
                     1936 => "00001100",
                     1937 => "01000111",
                     1938 => "00100100",
                     1939 => "00100011",
                     1940 => "11011100",
                     1941 => "00000001",
                     1942 => "10111010",
                     1943 => "11111111",
                     1944 => "00100001",
                     1945 => "11001101",
                     1946 => "00000101",
                     1947 => "00010110",
                     1948 => "00001010",
                     1949 => "00011011",
                     1950 => "00010010",
                     1951 => "00011000",
                     1952 => "00100010",
                     1953 => "00001100",
                     1954 => "00000111",
                     1955 => "00011101",
                     1956 => "00010010",
                     1957 => "00010110",
                     1958 => "00001110",
                     1959 => "00100100",
                     1960 => "00011110",
                     1961 => "00011001",
                     1962 => "11111111",
                     1963 => "00100001",
                     1964 => "11001101",
                     1965 => "00000101",
                     1966 => "00010110",
                     1967 => "00001010",
                     1968 => "00011011",
                     1969 => "00010010",
                     1970 => "00011000",
                     1971 => "00100010",
                     1972 => "00001011",
                     1973 => "00001001",
                     1974 => "00010000",
                     1975 => "00001010",
                     1976 => "00010110",
                     1977 => "00001110",
                     1978 => "00100100",
                     1979 => "00011000",
                     1980 => "00011111",
                     1981 => "00001110",
                     1982 => "00011011",
                     1983 => "11111111",
                     1984 => "00100101",
                     1985 => "10000100",
                     1986 => "00010101",
                     1987 => "00100000",
                     1988 => "00001110",
                     1989 => "00010101",
                     1990 => "00001100",
                     1991 => "00011000",
                     1992 => "00010110",
                     1993 => "00001110",
                     1994 => "00100100",
                     1995 => "00011101",
                     1996 => "00011000",
                     1997 => "00100100",
                     1998 => "00100000",
                     1999 => "00001010",
                     2000 => "00011011",
                     2001 => "00011001",
                     2002 => "00100100",
                     2003 => "00100011",
                     2004 => "00011000",
                     2005 => "00010111",
                     2006 => "00001110",
                     2007 => "00101011",
                     2008 => "00100110",
                     2009 => "00100101",
                     2010 => "00000001",
                     2011 => "00100100",
                     2012 => "00100110",
                     2013 => "00101101",
                     2014 => "00000001",
                     2015 => "00100100",
                     2016 => "00100110",
                     2017 => "00110101",
                     2018 => "00000001",
                     2019 => "00100100",
                     2020 => "00100111",
                     2021 => "11011001",
                     2022 => "01000110",
                     2023 => "10101010",
                     2024 => "00100111",
                     2025 => "11100001",
                     2026 => "01000101",
                     2027 => "10101010",
                     2028 => "11111111",
                     2029 => "00010101",
                     2030 => "00011110",
                     2031 => "00010010",
                     2032 => "00010000",
                     2033 => "00010010",
                     2034 => "00000100",
                     2035 => "00000011",
                     2036 => "00000010",
                     2037 => "00000000",
                     2038 => "00100100",
                     2039 => "00000101",
                     2040 => "00100100",
                     2041 => "00000000",
                     2042 => "00001000",
                     2043 => "00000111",
                     2044 => "00000110",
                     2045 => "00000000",
                     2046 => "00000000",
                     2047 => "00000000",
                     2048 => "00100111",
                     2049 => "00100111",
                     2050 => "01000110",
                     2051 => "01001110",
                     2052 => "01011001",
                     2053 => "01100001",
                     2054 => "01101110",
                     2055 => "01101110",
                     2056 => "01001000",
                     2057 => "00001010",
                     2058 => "10101000",
                     2059 => "11000000",
                     2060 => "00000100",
                     2061 => "10010000",
                     2062 => "00001100",
                     2063 => "11000000",
                     2064 => "00001000",
                     2065 => "10010000",
                     2066 => "00000010",
                     2067 => "10100000",
                     2068 => "00001000",
                     2069 => "10101101",
                     2070 => "01111010",
                     2071 => "00000111",
                     2072 => "11010000",
                     2073 => "00000001",
                     2074 => "11001000",
                     2075 => "10111110",
                     2076 => "11111110",
                     2077 => "10000111",
                     2078 => "10100000",
                     2079 => "00000000",
                     2080 => "10111101",
                     2081 => "01010010",
                     2082 => "10000111",
                     2083 => "11001001",
                     2084 => "11111111",
                     2085 => "11110000",
                     2086 => "00000111",
                     2087 => "10011001",
                     2088 => "00000001",
                     2089 => "00000011",
                     2090 => "11101000",
                     2091 => "11001000",
                     2092 => "11010000",
                     2093 => "11110010",
                     2094 => "10101001",
                     2095 => "00000000",
                     2096 => "10011001",
                     2097 => "00000001",
                     2098 => "00000011",
                     2099 => "01101000",
                     2100 => "10101010",
                     2101 => "11001001",
                     2102 => "00000100",
                     2103 => "10110000",
                     2104 => "01001001",
                     2105 => "11001010",
                     2106 => "11010000",
                     2107 => "00100011",
                     2108 => "10101101",
                     2109 => "01011010",
                     2110 => "00000111",
                     2111 => "00011000",
                     2112 => "01101001",
                     2113 => "00000001",
                     2114 => "11001001",
                     2115 => "00001010",
                     2116 => "10010000",
                     2117 => "00000111",
                     2118 => "11101001",
                     2119 => "00001010",
                     2120 => "10100000",
                     2121 => "10011111",
                     2122 => "10001100",
                     2123 => "00001000",
                     2124 => "00000011",
                     2125 => "10001101",
                     2126 => "00001001",
                     2127 => "00000011",
                     2128 => "10101100",
                     2129 => "01011111",
                     2130 => "00000111",
                     2131 => "11001000",
                     2132 => "10001100",
                     2133 => "00010100",
                     2134 => "00000011",
                     2135 => "10101100",
                     2136 => "01011100",
                     2137 => "00000111",
                     2138 => "11001000",
                     2139 => "10001100",
                     2140 => "00010110",
                     2141 => "00000011",
                     2142 => "01100000",
                     2143 => "10101101",
                     2144 => "01111010",
                     2145 => "00000111",
                     2146 => "11110000",
                     2147 => "00011101",
                     2148 => "10101101",
                     2149 => "01010011",
                     2150 => "00000111",
                     2151 => "11001010",
                     2152 => "11010000",
                     2153 => "00001001",
                     2154 => "10101100",
                     2155 => "01110000",
                     2156 => "00000111",
                     2157 => "11000000",
                     2158 => "00000011",
                     2159 => "11110000",
                     2160 => "00000010",
                     2161 => "01001001",
                     2162 => "00000001",
                     2163 => "01001010",
                     2164 => "10010000",
                     2165 => "00001011",
                     2166 => "10100000",
                     2167 => "00000100",
                     2168 => "10111001",
                     2169 => "11101101",
                     2170 => "10000111",
                     2171 => "10011001",
                     2172 => "00000100",
                     2173 => "00000011",
                     2174 => "10001000",
                     2175 => "00010000",
                     2176 => "11110111",
                     2177 => "01100000",
                     2178 => "11101001",
                     2179 => "00000100",
                     2180 => "00001010",
                     2181 => "00001010",
                     2182 => "10101010",
                     2183 => "10100000",
                     2184 => "00000000",
                     2185 => "10111101",
                     2186 => "11110010",
                     2187 => "10000111",
                     2188 => "10011001",
                     2189 => "00011100",
                     2190 => "00000011",
                     2191 => "11101000",
                     2192 => "11001000",
                     2193 => "11001000",
                     2194 => "11001000",
                     2195 => "11001000",
                     2196 => "11000000",
                     2197 => "00001100",
                     2198 => "10010000",
                     2199 => "11110001",
                     2200 => "10101001",
                     2201 => "00101100",
                     2202 => "01001100",
                     2203 => "00111111",
                     2204 => "10000110",
                     2205 => "10101101",
                     2206 => "10100000",
                     2207 => "00000111",
                     2208 => "11010000",
                     2209 => "00001011",
                     2210 => "00100000",
                     2211 => "00100000",
                     2212 => "10000010",
                     2213 => "10101001",
                     2214 => "00000111",
                     2215 => "10001101",
                     2216 => "10100000",
                     2217 => "00000111",
                     2218 => "11101110",
                     2219 => "00111100",
                     2220 => "00000111",
                     2221 => "01100000",
                     2222 => "10101101",
                     2223 => "00100110",
                     2224 => "00000111",
                     2225 => "00101001",
                     2226 => "00000001",
                     2227 => "10000101",
                     2228 => "00000101",
                     2229 => "10101100",
                     2230 => "01000000",
                     2231 => "00000011",
                     2232 => "10000100",
                     2233 => "00000000",
                     2234 => "10101101",
                     2235 => "00100001",
                     2236 => "00000111",
                     2237 => "10011001",
                     2238 => "01000010",
                     2239 => "00000011",
                     2240 => "10101101",
                     2241 => "00100000",
                     2242 => "00000111",
                     2243 => "10011001",
                     2244 => "01000001",
                     2245 => "00000011",
                     2246 => "10101001",
                     2247 => "10011010",
                     2248 => "10011001",
                     2249 => "01000011",
                     2250 => "00000011",
                     2251 => "10101001",
                     2252 => "00000000",
                     2253 => "10000101",
                     2254 => "00000100",
                     2255 => "10101010",
                     2256 => "10000110",
                     2257 => "00000001",
                     2258 => "10111101",
                     2259 => "10100001",
                     2260 => "00000110",
                     2261 => "00101001",
                     2262 => "11000000",
                     2263 => "10000101",
                     2264 => "00000011",
                     2265 => "00001010",
                     2266 => "00101010",
                     2267 => "00101010",
                     2268 => "10101000",
                     2269 => "10111001",
                     2270 => "00001000",
                     2271 => "10001011",
                     2272 => "10000101",
                     2273 => "00000110",
                     2274 => "10111001",
                     2275 => "00001100",
                     2276 => "10001011",
                     2277 => "10000101",
                     2278 => "00000111",
                     2279 => "10111101",
                     2280 => "10100001",
                     2281 => "00000110",
                     2282 => "00001010",
                     2283 => "00001010",
                     2284 => "10000101",
                     2285 => "00000010",
                     2286 => "10101101",
                     2287 => "00011111",
                     2288 => "00000111",
                     2289 => "00101001",
                     2290 => "00000001",
                     2291 => "01001001",
                     2292 => "00000001",
                     2293 => "00001010",
                     2294 => "01100101",
                     2295 => "00000010",
                     2296 => "10101000",
                     2297 => "10100110",
                     2298 => "00000000",
                     2299 => "10110001",
                     2300 => "00000110",
                     2301 => "10011101",
                     2302 => "01000100",
                     2303 => "00000011",
                     2304 => "11001000",
                     2305 => "10110001",
                     2306 => "00000110",
                     2307 => "10011101",
                     2308 => "01000101",
                     2309 => "00000011",
                     2310 => "10100100",
                     2311 => "00000100",
                     2312 => "10100101",
                     2313 => "00000101",
                     2314 => "11010000",
                     2315 => "00001110",
                     2316 => "10100101",
                     2317 => "00000001",
                     2318 => "01001010",
                     2319 => "10110000",
                     2320 => "00011001",
                     2321 => "00100110",
                     2322 => "00000011",
                     2323 => "00100110",
                     2324 => "00000011",
                     2325 => "00100110",
                     2326 => "00000011",
                     2327 => "01001100",
                     2328 => "00110000",
                     2329 => "10001001",
                     2330 => "10100101",
                     2331 => "00000001",
                     2332 => "01001010",
                     2333 => "10110000",
                     2334 => "00001111",
                     2335 => "01000110",
                     2336 => "00000011",
                     2337 => "01000110",
                     2338 => "00000011",
                     2339 => "01000110",
                     2340 => "00000011",
                     2341 => "01000110",
                     2342 => "00000011",
                     2343 => "01001100",
                     2344 => "00110000",
                     2345 => "10001001",
                     2346 => "01000110",
                     2347 => "00000011",
                     2348 => "01000110",
                     2349 => "00000011",
                     2350 => "11100110",
                     2351 => "00000100",
                     2352 => "10111001",
                     2353 => "11111001",
                     2354 => "00000011",
                     2355 => "00000101",
                     2356 => "00000011",
                     2357 => "10011001",
                     2358 => "11111001",
                     2359 => "00000011",
                     2360 => "11100110",
                     2361 => "00000000",
                     2362 => "11100110",
                     2363 => "00000000",
                     2364 => "10100110",
                     2365 => "00000001",
                     2366 => "11101000",
                     2367 => "11100000",
                     2368 => "00001101",
                     2369 => "10010000",
                     2370 => "10001101",
                     2371 => "10100100",
                     2372 => "00000000",
                     2373 => "11001000",
                     2374 => "11001000",
                     2375 => "11001000",
                     2376 => "10101001",
                     2377 => "00000000",
                     2378 => "10011001",
                     2379 => "01000001",
                     2380 => "00000011",
                     2381 => "10001100",
                     2382 => "01000000",
                     2383 => "00000011",
                     2384 => "11101110",
                     2385 => "00100001",
                     2386 => "00000111",
                     2387 => "10101101",
                     2388 => "00100001",
                     2389 => "00000111",
                     2390 => "00101001",
                     2391 => "00011111",
                     2392 => "11010000",
                     2393 => "00001101",
                     2394 => "10101001",
                     2395 => "10000000",
                     2396 => "10001101",
                     2397 => "00100001",
                     2398 => "00000111",
                     2399 => "10101101",
                     2400 => "00100000",
                     2401 => "00000111",
                     2402 => "01001001",
                     2403 => "00000100",
                     2404 => "10001101",
                     2405 => "00100000",
                     2406 => "00000111",
                     2407 => "01001100",
                     2408 => "10111101",
                     2409 => "10001001",
                     2410 => "10101101",
                     2411 => "00100001",
                     2412 => "00000111",
                     2413 => "00101001",
                     2414 => "00011111",
                     2415 => "00111000",
                     2416 => "11101001",
                     2417 => "00000100",
                     2418 => "00101001",
                     2419 => "00011111",
                     2420 => "10000101",
                     2421 => "00000001",
                     2422 => "10101101",
                     2423 => "00100000",
                     2424 => "00000111",
                     2425 => "10110000",
                     2426 => "00000010",
                     2427 => "01001001",
                     2428 => "00000100",
                     2429 => "00101001",
                     2430 => "00000100",
                     2431 => "00001001",
                     2432 => "00100011",
                     2433 => "10000101",
                     2434 => "00000000",
                     2435 => "10100101",
                     2436 => "00000001",
                     2437 => "01001010",
                     2438 => "01001010",
                     2439 => "01101001",
                     2440 => "11000000",
                     2441 => "10000101",
                     2442 => "00000001",
                     2443 => "10100010",
                     2444 => "00000000",
                     2445 => "10101100",
                     2446 => "01000000",
                     2447 => "00000011",
                     2448 => "10100101",
                     2449 => "00000000",
                     2450 => "10011001",
                     2451 => "01000001",
                     2452 => "00000011",
                     2453 => "10100101",
                     2454 => "00000001",
                     2455 => "00011000",
                     2456 => "01101001",
                     2457 => "00001000",
                     2458 => "10011001",
                     2459 => "01000010",
                     2460 => "00000011",
                     2461 => "10000101",
                     2462 => "00000001",
                     2463 => "10111101",
                     2464 => "11111001",
                     2465 => "00000011",
                     2466 => "10011001",
                     2467 => "01000100",
                     2468 => "00000011",
                     2469 => "10101001",
                     2470 => "00000001",
                     2471 => "10011001",
                     2472 => "01000011",
                     2473 => "00000011",
                     2474 => "01001010",
                     2475 => "10011101",
                     2476 => "11111001",
                     2477 => "00000011",
                     2478 => "11001000",
                     2479 => "11001000",
                     2480 => "11001000",
                     2481 => "11001000",
                     2482 => "11101000",
                     2483 => "11100000",
                     2484 => "00000111",
                     2485 => "10010000",
                     2486 => "11011001",
                     2487 => "10011001",
                     2488 => "01000001",
                     2489 => "00000011",
                     2490 => "10001100",
                     2491 => "01000000",
                     2492 => "00000011",
                     2493 => "10101001",
                     2494 => "00000110",
                     2495 => "10001101",
                     2496 => "01110011",
                     2497 => "00000111",
                     2498 => "01100000",
                     2499 => "00100111",
                     2500 => "00100111",
                     2501 => "00100111",
                     2502 => "00010111",
                     2503 => "00000111",
                     2504 => "00010111",
                     2505 => "00111111",
                     2506 => "00001100",
                     2507 => "00000100",
                     2508 => "11111111",
                     2509 => "11111111",
                     2510 => "11111111",
                     2511 => "11111111",
                     2512 => "00000000",
                     2513 => "00001111",
                     2514 => "00000111",
                     2515 => "00010010",
                     2516 => "00001111",
                     2517 => "00001111",
                     2518 => "00000111",
                     2519 => "00010111",
                     2520 => "00001111",
                     2521 => "00001111",
                     2522 => "00000111",
                     2523 => "00010111",
                     2524 => "00011100",
                     2525 => "00001111",
                     2526 => "00000111",
                     2527 => "00010111",
                     2528 => "00000000",
                     2529 => "10100101",
                     2530 => "00001001",
                     2531 => "00101001",
                     2532 => "00000111",
                     2533 => "11010000",
                     2534 => "01010001",
                     2535 => "10101110",
                     2536 => "00000000",
                     2537 => "00000011",
                     2538 => "11100000",
                     2539 => "00110001",
                     2540 => "10110000",
                     2541 => "01001010",
                     2542 => "10101000",
                     2543 => "10111001",
                     2544 => "11001001",
                     2545 => "10001001",
                     2546 => "10011101",
                     2547 => "00000001",
                     2548 => "00000011",
                     2549 => "11101000",
                     2550 => "11001000",
                     2551 => "11000000",
                     2552 => "00001000",
                     2553 => "10010000",
                     2554 => "11110100",
                     2555 => "10101110",
                     2556 => "00000000",
                     2557 => "00000011",
                     2558 => "10101001",
                     2559 => "00000011",
                     2560 => "10000101",
                     2561 => "00000000",
                     2562 => "10101101",
                     2563 => "01001110",
                     2564 => "00000111",
                     2565 => "00001010",
                     2566 => "00001010",
                     2567 => "10101000",
                     2568 => "10111001",
                     2569 => "11010001",
                     2570 => "10001001",
                     2571 => "10011101",
                     2572 => "00000100",
                     2573 => "00000011",
                     2574 => "11001000",
                     2575 => "11101000",
                     2576 => "11000110",
                     2577 => "00000000",
                     2578 => "00010000",
                     2579 => "11110100",
                     2580 => "10101110",
                     2581 => "00000000",
                     2582 => "00000011",
                     2583 => "10101100",
                     2584 => "11010100",
                     2585 => "00000110",
                     2586 => "10111001",
                     2587 => "11000011",
                     2588 => "10001001",
                     2589 => "10011101",
                     2590 => "00000101",
                     2591 => "00000011",
                     2592 => "10101101",
                     2593 => "00000000",
                     2594 => "00000011",
                     2595 => "00011000",
                     2596 => "01101001",
                     2597 => "00000111",
                     2598 => "10001101",
                     2599 => "00000000",
                     2600 => "00000011",
                     2601 => "11101110",
                     2602 => "11010100",
                     2603 => "00000110",
                     2604 => "10101101",
                     2605 => "11010100",
                     2606 => "00000110",
                     2607 => "11001001",
                     2608 => "00000110",
                     2609 => "10010000",
                     2610 => "00000101",
                     2611 => "10101001",
                     2612 => "00000000",
                     2613 => "10001101",
                     2614 => "11010100",
                     2615 => "00000110",
                     2616 => "01100000",
                     2617 => "01000101",
                     2618 => "01000101",
                     2619 => "01000111",
                     2620 => "01000111",
                     2621 => "01000111",
                     2622 => "01000111",
                     2623 => "01000111",
                     2624 => "01000111",
                     2625 => "01010111",
                     2626 => "01011000",
                     2627 => "01011001",
                     2628 => "01011010",
                     2629 => "00100100",
                     2630 => "00100100",
                     2631 => "00100100",
                     2632 => "00100100",
                     2633 => "00100110",
                     2634 => "00100110",
                     2635 => "00100110",
                     2636 => "00100110",
                     2637 => "10100000",
                     2638 => "01000001",
                     2639 => "10101001",
                     2640 => "00000011",
                     2641 => "10101110",
                     2642 => "01001110",
                     2643 => "00000111",
                     2644 => "11010000",
                     2645 => "00000010",
                     2646 => "10101001",
                     2647 => "00000100",
                     2648 => "00100000",
                     2649 => "10010111",
                     2650 => "10001010",
                     2651 => "10101001",
                     2652 => "00000110",
                     2653 => "10001101",
                     2654 => "01110011",
                     2655 => "00000111",
                     2656 => "01100000",
                     2657 => "00100000",
                     2658 => "01101101",
                     2659 => "10001010",
                     2660 => "11101110",
                     2661 => "11110000",
                     2662 => "00000011",
                     2663 => "11011110",
                     2664 => "11101100",
                     2665 => "00000011",
                     2666 => "01100000",
                     2667 => "10101001",
                     2668 => "00000000",
                     2669 => "10100000",
                     2670 => "00000011",
                     2671 => "11001001",
                     2672 => "00000000",
                     2673 => "11110000",
                     2674 => "00010100",
                     2675 => "10100000",
                     2676 => "00000000",
                     2677 => "11001001",
                     2678 => "01011000",
                     2679 => "11110000",
                     2680 => "00001110",
                     2681 => "11001001",
                     2682 => "01010001",
                     2683 => "11110000",
                     2684 => "00001010",
                     2685 => "11001000",
                     2686 => "11001001",
                     2687 => "01011101",
                     2688 => "11110000",
                     2689 => "00000101",
                     2690 => "11001001",
                     2691 => "01010010",
                     2692 => "11110000",
                     2693 => "00000001",
                     2694 => "11001000",
                     2695 => "10011000",
                     2696 => "10101100",
                     2697 => "00000000",
                     2698 => "00000011",
                     2699 => "11001000",
                     2700 => "00100000",
                     2701 => "10010111",
                     2702 => "10001010",
                     2703 => "10001000",
                     2704 => "10011000",
                     2705 => "00011000",
                     2706 => "01101001",
                     2707 => "00001010",
                     2708 => "01001100",
                     2709 => "00111111",
                     2710 => "10000110",
                     2711 => "10000110",
                     2712 => "00000000",
                     2713 => "10000100",
                     2714 => "00000001",
                     2715 => "00001010",
                     2716 => "00001010",
                     2717 => "10101010",
                     2718 => "10100000",
                     2719 => "00100000",
                     2720 => "10100101",
                     2721 => "00000110",
                     2722 => "11001001",
                     2723 => "11010000",
                     2724 => "10010000",
                     2725 => "00000010",
                     2726 => "10100000",
                     2727 => "00100100",
                     2728 => "10000100",
                     2729 => "00000011",
                     2730 => "00101001",
                     2731 => "00001111",
                     2732 => "00001010",
                     2733 => "10000101",
                     2734 => "00000100",
                     2735 => "10101001",
                     2736 => "00000000",
                     2737 => "10000101",
                     2738 => "00000101",
                     2739 => "10100101",
                     2740 => "00000010",
                     2741 => "00011000",
                     2742 => "01101001",
                     2743 => "00100000",
                     2744 => "00001010",
                     2745 => "00100110",
                     2746 => "00000101",
                     2747 => "00001010",
                     2748 => "00100110",
                     2749 => "00000101",
                     2750 => "01100101",
                     2751 => "00000100",
                     2752 => "10000101",
                     2753 => "00000100",
                     2754 => "10100101",
                     2755 => "00000101",
                     2756 => "01101001",
                     2757 => "00000000",
                     2758 => "00011000",
                     2759 => "01100101",
                     2760 => "00000011",
                     2761 => "10000101",
                     2762 => "00000101",
                     2763 => "10100100",
                     2764 => "00000001",
                     2765 => "10111101",
                     2766 => "00111001",
                     2767 => "10001010",
                     2768 => "10011001",
                     2769 => "00000011",
                     2770 => "00000011",
                     2771 => "10111101",
                     2772 => "00111010",
                     2773 => "10001010",
                     2774 => "10011001",
                     2775 => "00000100",
                     2776 => "00000011",
                     2777 => "10111101",
                     2778 => "00111011",
                     2779 => "10001010",
                     2780 => "10011001",
                     2781 => "00001000",
                     2782 => "00000011",
                     2783 => "10111101",
                     2784 => "00111100",
                     2785 => "10001010",
                     2786 => "10011001",
                     2787 => "00001001",
                     2788 => "00000011",
                     2789 => "10100101",
                     2790 => "00000100",
                     2791 => "10011001",
                     2792 => "00000001",
                     2793 => "00000011",
                     2794 => "00011000",
                     2795 => "01101001",
                     2796 => "00100000",
                     2797 => "10011001",
                     2798 => "00000110",
                     2799 => "00000011",
                     2800 => "10100101",
                     2801 => "00000101",
                     2802 => "10011001",
                     2803 => "00000000",
                     2804 => "00000011",
                     2805 => "10011001",
                     2806 => "00000101",
                     2807 => "00000011",
                     2808 => "10101001",
                     2809 => "00000010",
                     2810 => "10011001",
                     2811 => "00000010",
                     2812 => "00000011",
                     2813 => "10011001",
                     2814 => "00000111",
                     2815 => "00000011",
                     2816 => "10101001",
                     2817 => "00000000",
                     2818 => "10011001",
                     2819 => "00001010",
                     2820 => "00000011",
                     2821 => "10100110",
                     2822 => "00000000",
                     2823 => "01100000",
                     2824 => "00010000",
                     2825 => "10101100",
                     2826 => "01100100",
                     2827 => "10001100",
                     2828 => "10001011",
                     2829 => "10001011",
                     2830 => "10001100",
                     2831 => "10001100",
                     2832 => "00100100",
                     2833 => "00100100",
                     2834 => "00100100",
                     2835 => "00100100",
                     2836 => "00100111",
                     2837 => "00100111",
                     2838 => "00100111",
                     2839 => "00100111",
                     2840 => "00100100",
                     2841 => "00100100",
                     2842 => "00100100",
                     2843 => "00110101",
                     2844 => "00110110",
                     2845 => "00100101",
                     2846 => "00110111",
                     2847 => "00100101",
                     2848 => "00100100",
                     2849 => "00111000",
                     2850 => "00100100",
                     2851 => "00100100",
                     2852 => "00100100",
                     2853 => "00110000",
                     2854 => "00110000",
                     2855 => "00100110",
                     2856 => "00100110",
                     2857 => "00100110",
                     2858 => "00110100",
                     2859 => "00100110",
                     2860 => "00100100",
                     2861 => "00110001",
                     2862 => "00100100",
                     2863 => "00110010",
                     2864 => "00110011",
                     2865 => "00100110",
                     2866 => "00100100",
                     2867 => "00110011",
                     2868 => "00110100",
                     2869 => "00100110",
                     2870 => "00100110",
                     2871 => "00100110",
                     2872 => "00100110",
                     2873 => "00100110",
                     2874 => "00100110",
                     2875 => "00100110",
                     2876 => "00100100",
                     2877 => "11000000",
                     2878 => "00100100",
                     2879 => "11000000",
                     2880 => "00100100",
                     2881 => "01111111",
                     2882 => "01111111",
                     2883 => "00100100",
                     2884 => "10111000",
                     2885 => "10111010",
                     2886 => "10111001",
                     2887 => "10111011",
                     2888 => "10111000",
                     2889 => "10111100",
                     2890 => "10111001",
                     2891 => "10111101",
                     2892 => "10111010",
                     2893 => "10111100",
                     2894 => "10111011",
                     2895 => "10111101",
                     2896 => "01100000",
                     2897 => "01100100",
                     2898 => "01100001",
                     2899 => "01100101",
                     2900 => "01100010",
                     2901 => "01100110",
                     2902 => "01100011",
                     2903 => "01100111",
                     2904 => "01100000",
                     2905 => "01100100",
                     2906 => "01100001",
                     2907 => "01100101",
                     2908 => "01100010",
                     2909 => "01100110",
                     2910 => "01100011",
                     2911 => "01100111",
                     2912 => "01101000",
                     2913 => "01101000",
                     2914 => "01101001",
                     2915 => "01101001",
                     2916 => "00100110",
                     2917 => "00100110",
                     2918 => "01101010",
                     2919 => "01101010",
                     2920 => "01001011",
                     2921 => "01001100",
                     2922 => "01001101",
                     2923 => "01001110",
                     2924 => "01001101",
                     2925 => "01001111",
                     2926 => "01001101",
                     2927 => "01001111",
                     2928 => "01001101",
                     2929 => "01001110",
                     2930 => "01010000",
                     2931 => "01010001",
                     2932 => "01101011",
                     2933 => "01110000",
                     2934 => "00101100",
                     2935 => "00101101",
                     2936 => "01101100",
                     2937 => "01110001",
                     2938 => "01101101",
                     2939 => "01110010",
                     2940 => "01101110",
                     2941 => "01110011",
                     2942 => "01101111",
                     2943 => "01110100",
                     2944 => "10000110",
                     2945 => "10001010",
                     2946 => "10000111",
                     2947 => "10001011",
                     2948 => "10001000",
                     2949 => "10001100",
                     2950 => "10001000",
                     2951 => "10001100",
                     2952 => "10001001",
                     2953 => "10001101",
                     2954 => "01101001",
                     2955 => "01101001",
                     2956 => "10001110",
                     2957 => "10010001",
                     2958 => "10001111",
                     2959 => "10010010",
                     2960 => "00100110",
                     2961 => "10010011",
                     2962 => "00100110",
                     2963 => "10010011",
                     2964 => "10010000",
                     2965 => "10010100",
                     2966 => "01101001",
                     2967 => "01101001",
                     2968 => "10100100",
                     2969 => "11101001",
                     2970 => "11101010",
                     2971 => "11101011",
                     2972 => "00100100",
                     2973 => "00100100",
                     2974 => "00100100",
                     2975 => "00100100",
                     2976 => "00100100",
                     2977 => "00101111",
                     2978 => "00100100",
                     2979 => "00111101",
                     2980 => "10100010",
                     2981 => "10100010",
                     2982 => "10100011",
                     2983 => "10100011",
                     2984 => "00100100",
                     2985 => "00100100",
                     2986 => "00100100",
                     2987 => "00100100",
                     2988 => "10100010",
                     2989 => "10100010",
                     2990 => "10100011",
                     2991 => "10100011",
                     2992 => "10011001",
                     2993 => "00100100",
                     2994 => "10011001",
                     2995 => "00100100",
                     2996 => "00100100",
                     2997 => "10100010",
                     2998 => "00111110",
                     2999 => "00111111",
                     3000 => "01011011",
                     3001 => "01011100",
                     3002 => "00100100",
                     3003 => "10100011",
                     3004 => "00100100",
                     3005 => "00100100",
                     3006 => "00100100",
                     3007 => "00100100",
                     3008 => "10011101",
                     3009 => "01000111",
                     3010 => "10011110",
                     3011 => "01000111",
                     3012 => "01000111",
                     3013 => "01000111",
                     3014 => "00100111",
                     3015 => "00100111",
                     3016 => "01000111",
                     3017 => "01000111",
                     3018 => "01000111",
                     3019 => "01000111",
                     3020 => "00100111",
                     3021 => "00100111",
                     3022 => "01000111",
                     3023 => "01000111",
                     3024 => "10101001",
                     3025 => "01000111",
                     3026 => "10101010",
                     3027 => "01000111",
                     3028 => "10011011",
                     3029 => "00100111",
                     3030 => "10011100",
                     3031 => "00100111",
                     3032 => "00100111",
                     3033 => "00100111",
                     3034 => "00100111",
                     3035 => "00100111",
                     3036 => "01010010",
                     3037 => "01010010",
                     3038 => "01010010",
                     3039 => "01010010",
                     3040 => "10000000",
                     3041 => "10100000",
                     3042 => "10000001",
                     3043 => "10100001",
                     3044 => "10111110",
                     3045 => "10111110",
                     3046 => "10111111",
                     3047 => "10111111",
                     3048 => "01110101",
                     3049 => "10111010",
                     3050 => "01110110",
                     3051 => "10111011",
                     3052 => "10111010",
                     3053 => "10111010",
                     3054 => "10111011",
                     3055 => "10111011",
                     3056 => "01000101",
                     3057 => "01000111",
                     3058 => "01000101",
                     3059 => "01000111",
                     3060 => "01000111",
                     3061 => "01000111",
                     3062 => "01000111",
                     3063 => "01000111",
                     3064 => "01000101",
                     3065 => "01000111",
                     3066 => "01000101",
                     3067 => "01000111",
                     3068 => "10110100",
                     3069 => "10110110",
                     3070 => "10110101",
                     3071 => "10110111",
                     3072 => "01000101",
                     3073 => "01000111",
                     3074 => "01000101",
                     3075 => "01000111",
                     3076 => "01000101",
                     3077 => "01000111",
                     3078 => "01000101",
                     3079 => "01000111",
                     3080 => "01000101",
                     3081 => "01000111",
                     3082 => "01000101",
                     3083 => "01000111",
                     3084 => "01000101",
                     3085 => "01000111",
                     3086 => "01000101",
                     3087 => "01000111",
                     3088 => "01000101",
                     3089 => "01000111",
                     3090 => "01000101",
                     3091 => "01000111",
                     3092 => "01000111",
                     3093 => "01000111",
                     3094 => "01000111",
                     3095 => "01000111",
                     3096 => "01000111",
                     3097 => "01000111",
                     3098 => "01000111",
                     3099 => "01000111",
                     3100 => "01000111",
                     3101 => "01000111",
                     3102 => "01000111",
                     3103 => "01000111",
                     3104 => "01000111",
                     3105 => "01000111",
                     3106 => "01000111",
                     3107 => "01000111",
                     3108 => "01000111",
                     3109 => "01000111",
                     3110 => "01000111",
                     3111 => "01000111",
                     3112 => "00100100",
                     3113 => "00100100",
                     3114 => "00100100",
                     3115 => "00100100",
                     3116 => "00100100",
                     3117 => "00100100",
                     3118 => "00100100",
                     3119 => "00100100",
                     3120 => "10101011",
                     3121 => "10101100",
                     3122 => "10101101",
                     3123 => "10101110",
                     3124 => "01011101",
                     3125 => "01011110",
                     3126 => "01011101",
                     3127 => "01011110",
                     3128 => "11000001",
                     3129 => "00100100",
                     3130 => "11000001",
                     3131 => "00100100",
                     3132 => "11000110",
                     3133 => "11001000",
                     3134 => "11000111",
                     3135 => "11001001",
                     3136 => "11001010",
                     3137 => "11001100",
                     3138 => "11001011",
                     3139 => "11001101",
                     3140 => "00101010",
                     3141 => "00101010",
                     3142 => "01000000",
                     3143 => "01000000",
                     3144 => "00100100",
                     3145 => "00100100",
                     3146 => "00100100",
                     3147 => "00100100",
                     3148 => "00100100",
                     3149 => "01000111",
                     3150 => "00100100",
                     3151 => "01000111",
                     3152 => "10000010",
                     3153 => "10000011",
                     3154 => "10000100",
                     3155 => "10000101",
                     3156 => "00100100",
                     3157 => "01000111",
                     3158 => "00100100",
                     3159 => "01000111",
                     3160 => "10000110",
                     3161 => "10001010",
                     3162 => "10000111",
                     3163 => "10001011",
                     3164 => "10001110",
                     3165 => "10010001",
                     3166 => "10001111",
                     3167 => "10010010",
                     3168 => "00100100",
                     3169 => "00101111",
                     3170 => "00100100",
                     3171 => "00111101",
                     3172 => "00100100",
                     3173 => "00100100",
                     3174 => "00100100",
                     3175 => "00110101",
                     3176 => "00110110",
                     3177 => "00100101",
                     3178 => "00110111",
                     3179 => "00100101",
                     3180 => "00100100",
                     3181 => "00111000",
                     3182 => "00100100",
                     3183 => "00100100",
                     3184 => "00100100",
                     3185 => "00100100",
                     3186 => "00111001",
                     3187 => "00100100",
                     3188 => "00111010",
                     3189 => "00100100",
                     3190 => "00111011",
                     3191 => "00100100",
                     3192 => "00111100",
                     3193 => "00100100",
                     3194 => "00100100",
                     3195 => "00100100",
                     3196 => "01000001",
                     3197 => "00100110",
                     3198 => "01000001",
                     3199 => "00100110",
                     3200 => "00100110",
                     3201 => "00100110",
                     3202 => "00100110",
                     3203 => "00100110",
                     3204 => "10110000",
                     3205 => "10110001",
                     3206 => "10110010",
                     3207 => "10110011",
                     3208 => "01110111",
                     3209 => "01111001",
                     3210 => "01110111",
                     3211 => "01111001",
                     3212 => "01010011",
                     3213 => "01010101",
                     3214 => "01010100",
                     3215 => "01010110",
                     3216 => "01010011",
                     3217 => "01010101",
                     3218 => "01010100",
                     3219 => "01010110",
                     3220 => "10100101",
                     3221 => "10100111",
                     3222 => "10100110",
                     3223 => "10101000",
                     3224 => "11000010",
                     3225 => "11000100",
                     3226 => "11000011",
                     3227 => "11000101",
                     3228 => "01010111",
                     3229 => "01011001",
                     3230 => "01011000",
                     3231 => "01011010",
                     3232 => "01111011",
                     3233 => "01111101",
                     3234 => "01111100",
                     3235 => "01111110",
                     3236 => "00111111",
                     3237 => "00000000",
                     3238 => "00100000",
                     3239 => "00001111",
                     3240 => "00010101",
                     3241 => "00010010",
                     3242 => "00100101",
                     3243 => "00001111",
                     3244 => "00111010",
                     3245 => "00011010",
                     3246 => "00001111",
                     3247 => "00001111",
                     3248 => "00110000",
                     3249 => "00010010",
                     3250 => "00001111",
                     3251 => "00001111",
                     3252 => "00100111",
                     3253 => "00010010",
                     3254 => "00001111",
                     3255 => "00100010",
                     3256 => "00010110",
                     3257 => "00100111",
                     3258 => "00011000",
                     3259 => "00001111",
                     3260 => "00010000",
                     3261 => "00110000",
                     3262 => "00100111",
                     3263 => "00001111",
                     3264 => "00010110",
                     3265 => "00110000",
                     3266 => "00100111",
                     3267 => "00001111",
                     3268 => "00001111",
                     3269 => "00110000",
                     3270 => "00010000",
                     3271 => "00000000",
                     3272 => "00111111",
                     3273 => "00000000",
                     3274 => "00100000",
                     3275 => "00001111",
                     3276 => "00101001",
                     3277 => "00011010",
                     3278 => "00001111",
                     3279 => "00001111",
                     3280 => "00110110",
                     3281 => "00010111",
                     3282 => "00001111",
                     3283 => "00001111",
                     3284 => "00110000",
                     3285 => "00100001",
                     3286 => "00001111",
                     3287 => "00001111",
                     3288 => "00100111",
                     3289 => "00010111",
                     3290 => "00001111",
                     3291 => "00001111",
                     3292 => "00010110",
                     3293 => "00100111",
                     3294 => "00011000",
                     3295 => "00001111",
                     3296 => "00011010",
                     3297 => "00110000",
                     3298 => "00100111",
                     3299 => "00001111",
                     3300 => "00010110",
                     3301 => "00110000",
                     3302 => "00100111",
                     3303 => "00001111",
                     3304 => "00001111",
                     3305 => "00110110",
                     3306 => "00010111",
                     3307 => "00000000",
                     3308 => "00111111",
                     3309 => "00000000",
                     3310 => "00100000",
                     3311 => "00001111",
                     3312 => "00101001",
                     3313 => "00011010",
                     3314 => "00001001",
                     3315 => "00001111",
                     3316 => "00111100",
                     3317 => "00011100",
                     3318 => "00001111",
                     3319 => "00001111",
                     3320 => "00110000",
                     3321 => "00100001",
                     3322 => "00011100",
                     3323 => "00001111",
                     3324 => "00100111",
                     3325 => "00010111",
                     3326 => "00011100",
                     3327 => "00001111",
                     3328 => "00010110",
                     3329 => "00100111",
                     3330 => "00011000",
                     3331 => "00001111",
                     3332 => "00011100",
                     3333 => "00110110",
                     3334 => "00010111",
                     3335 => "00001111",
                     3336 => "00010110",
                     3337 => "00110000",
                     3338 => "00100111",
                     3339 => "00001111",
                     3340 => "00001100",
                     3341 => "00111100",
                     3342 => "00011100",
                     3343 => "00000000",
                     3344 => "00111111",
                     3345 => "00000000",
                     3346 => "00100000",
                     3347 => "00001111",
                     3348 => "00110000",
                     3349 => "00010000",
                     3350 => "00000000",
                     3351 => "00001111",
                     3352 => "00110000",
                     3353 => "00010000",
                     3354 => "00000000",
                     3355 => "00001111",
                     3356 => "00110000",
                     3357 => "00010110",
                     3358 => "00000000",
                     3359 => "00001111",
                     3360 => "00100111",
                     3361 => "00010111",
                     3362 => "00000000",
                     3363 => "00001111",
                     3364 => "00010110",
                     3365 => "00100111",
                     3366 => "00011000",
                     3367 => "00001111",
                     3368 => "00011100",
                     3369 => "00110110",
                     3370 => "00010111",
                     3371 => "00001111",
                     3372 => "00010110",
                     3373 => "00110000",
                     3374 => "00100111",
                     3375 => "00001111",
                     3376 => "00000000",
                     3377 => "00110000",
                     3378 => "00010000",
                     3379 => "00000000",
                     3380 => "00111111",
                     3381 => "00000000",
                     3382 => "00000100",
                     3383 => "00100010",
                     3384 => "00110000",
                     3385 => "00000000",
                     3386 => "00010000",
                     3387 => "00000000",
                     3388 => "00111111",
                     3389 => "00000000",
                     3390 => "00000100",
                     3391 => "00001111",
                     3392 => "00110000",
                     3393 => "00000000",
                     3394 => "00010000",
                     3395 => "00000000",
                     3396 => "00111111",
                     3397 => "00000000",
                     3398 => "00000100",
                     3399 => "00100010",
                     3400 => "00100111",
                     3401 => "00010110",
                     3402 => "00001111",
                     3403 => "00000000",
                     3404 => "00111111",
                     3405 => "00010100",
                     3406 => "00000100",
                     3407 => "00001111",
                     3408 => "00011010",
                     3409 => "00110000",
                     3410 => "00100111",
                     3411 => "00000000",
                     3412 => "00100101",
                     3413 => "01001000",
                     3414 => "00010000",
                     3415 => "00011101",
                     3416 => "00010001",
                     3417 => "00001010",
                     3418 => "00010111",
                     3419 => "00010100",
                     3420 => "00100100",
                     3421 => "00100010",
                     3422 => "00011000",
                     3423 => "00011110",
                     3424 => "00100100",
                     3425 => "00010110",
                     3426 => "00001010",
                     3427 => "00011011",
                     3428 => "00010010",
                     3429 => "00011000",
                     3430 => "00101011",
                     3431 => "00000000",
                     3432 => "00100101",
                     3433 => "01001000",
                     3434 => "00010000",
                     3435 => "00011101",
                     3436 => "00010001",
                     3437 => "00001010",
                     3438 => "00010111",
                     3439 => "00010100",
                     3440 => "00100100",
                     3441 => "00100010",
                     3442 => "00011000",
                     3443 => "00011110",
                     3444 => "00100100",
                     3445 => "00010101",
                     3446 => "00011110",
                     3447 => "00010010",
                     3448 => "00010000",
                     3449 => "00010010",
                     3450 => "00101011",
                     3451 => "00000000",
                     3452 => "00100101",
                     3453 => "11000101",
                     3454 => "00010110",
                     3455 => "00001011",
                     3456 => "00011110",
                     3457 => "00011101",
                     3458 => "00100100",
                     3459 => "00011000",
                     3460 => "00011110",
                     3461 => "00011011",
                     3462 => "00100100",
                     3463 => "00011001",
                     3464 => "00011011",
                     3465 => "00010010",
                     3466 => "00010111",
                     3467 => "00001100",
                     3468 => "00001110",
                     3469 => "00011100",
                     3470 => "00011100",
                     3471 => "00100100",
                     3472 => "00010010",
                     3473 => "00011100",
                     3474 => "00100100",
                     3475 => "00010010",
                     3476 => "00010111",
                     3477 => "00100110",
                     3478 => "00000101",
                     3479 => "00001111",
                     3480 => "00001010",
                     3481 => "00010111",
                     3482 => "00011000",
                     3483 => "00011101",
                     3484 => "00010001",
                     3485 => "00001110",
                     3486 => "00011011",
                     3487 => "00100100",
                     3488 => "00001100",
                     3489 => "00001010",
                     3490 => "00011100",
                     3491 => "00011101",
                     3492 => "00010101",
                     3493 => "00001110",
                     3494 => "00101011",
                     3495 => "00000000",
                     3496 => "00100101",
                     3497 => "10100111",
                     3498 => "00010011",
                     3499 => "00100010",
                     3500 => "00011000",
                     3501 => "00011110",
                     3502 => "00011011",
                     3503 => "00100100",
                     3504 => "00011010",
                     3505 => "00011110",
                     3506 => "00001110",
                     3507 => "00011100",
                     3508 => "00011101",
                     3509 => "00100100",
                     3510 => "00010010",
                     3511 => "00011100",
                     3512 => "00100100",
                     3513 => "00011000",
                     3514 => "00011111",
                     3515 => "00001110",
                     3516 => "00011011",
                     3517 => "10101111",
                     3518 => "00000000",
                     3519 => "00100101",
                     3520 => "11100011",
                     3521 => "00011011",
                     3522 => "00100000",
                     3523 => "00001110",
                     3524 => "00100100",
                     3525 => "00011001",
                     3526 => "00011011",
                     3527 => "00001110",
                     3528 => "00011100",
                     3529 => "00001110",
                     3530 => "00010111",
                     3531 => "00011101",
                     3532 => "00100100",
                     3533 => "00100010",
                     3534 => "00011000",
                     3535 => "00011110",
                     3536 => "00100100",
                     3537 => "00001010",
                     3538 => "00100100",
                     3539 => "00010111",
                     3540 => "00001110",
                     3541 => "00100000",
                     3542 => "00100100",
                     3543 => "00011010",
                     3544 => "00011110",
                     3545 => "00001110",
                     3546 => "00011100",
                     3547 => "00011101",
                     3548 => "10101111",
                     3549 => "00000000",
                     3550 => "00100110",
                     3551 => "01001010",
                     3552 => "00001101",
                     3553 => "00011001",
                     3554 => "00011110",
                     3555 => "00011100",
                     3556 => "00010001",
                     3557 => "00100100",
                     3558 => "00001011",
                     3559 => "00011110",
                     3560 => "00011101",
                     3561 => "00011101",
                     3562 => "00011000",
                     3563 => "00010111",
                     3564 => "00100100",
                     3565 => "00001011",
                     3566 => "00000000",
                     3567 => "00100110",
                     3568 => "10001000",
                     3569 => "00010001",
                     3570 => "00011101",
                     3571 => "00011000",
                     3572 => "00100100",
                     3573 => "00011100",
                     3574 => "00001110",
                     3575 => "00010101",
                     3576 => "00001110",
                     3577 => "00001100",
                     3578 => "00011101",
                     3579 => "00100100",
                     3580 => "00001010",
                     3581 => "00100100",
                     3582 => "00100000",
                     3583 => "00011000",
                     3584 => "00011011",
                     3585 => "00010101",
                     3586 => "00001101",
                     3587 => "00000000",
                     3588 => "00001010",
                     3589 => "10101000",
                     3590 => "01101000",
                     3591 => "10000101",
                     3592 => "00000100",
                     3593 => "01101000",
                     3594 => "10000101",
                     3595 => "00000101",
                     3596 => "11001000",
                     3597 => "10110001",
                     3598 => "00000100",
                     3599 => "10000101",
                     3600 => "00000110",
                     3601 => "11001000",
                     3602 => "10110001",
                     3603 => "00000100",
                     3604 => "10000101",
                     3605 => "00000111",
                     3606 => "01101100",
                     3607 => "00000110",
                     3608 => "00000000",
                     3609 => "10101101",
                     3610 => "00000010",
                     3611 => "00100000",
                     3612 => "10101101",
                     3613 => "01111000",
                     3614 => "00000111",
                     3615 => "00001001",
                     3616 => "00010000",
                     3617 => "00101001",
                     3618 => "11110000",
                     3619 => "00100000",
                     3620 => "11101101",
                     3621 => "10001110",
                     3622 => "10101001",
                     3623 => "00100100",
                     3624 => "00100000",
                     3625 => "00101101",
                     3626 => "10001110",
                     3627 => "10101001",
                     3628 => "00100000",
                     3629 => "10001101",
                     3630 => "00000110",
                     3631 => "00100000",
                     3632 => "10101001",
                     3633 => "00000000",
                     3634 => "10001101",
                     3635 => "00000110",
                     3636 => "00100000",
                     3637 => "10100010",
                     3638 => "00000100",
                     3639 => "10100000",
                     3640 => "11000000",
                     3641 => "10101001",
                     3642 => "00100100",
                     3643 => "10001101",
                     3644 => "00000111",
                     3645 => "00100000",
                     3646 => "10001000",
                     3647 => "11010000",
                     3648 => "11111010",
                     3649 => "11001010",
                     3650 => "11010000",
                     3651 => "11110111",
                     3652 => "10100000",
                     3653 => "01000000",
                     3654 => "10001010",
                     3655 => "10001101",
                     3656 => "00000000",
                     3657 => "00000011",
                     3658 => "10001101",
                     3659 => "00000001",
                     3660 => "00000011",
                     3661 => "10001101",
                     3662 => "00000111",
                     3663 => "00100000",
                     3664 => "10001000",
                     3665 => "11010000",
                     3666 => "11111010",
                     3667 => "10001101",
                     3668 => "00111111",
                     3669 => "00000111",
                     3670 => "10001101",
                     3671 => "01000000",
                     3672 => "00000111",
                     3673 => "01001100",
                     3674 => "11100110",
                     3675 => "10001110",
                     3676 => "10101001",
                     3677 => "00000001",
                     3678 => "10001101",
                     3679 => "00010110",
                     3680 => "01000000",
                     3681 => "01001010",
                     3682 => "10101010",
                     3683 => "10001101",
                     3684 => "00010110",
                     3685 => "01000000",
                     3686 => "00100000",
                     3687 => "01101010",
                     3688 => "10001110",
                     3689 => "11101000",
                     3690 => "10100000",
                     3691 => "00001000",
                     3692 => "01001000",
                     3693 => "10111101",
                     3694 => "00010110",
                     3695 => "01000000",
                     3696 => "10000101",
                     3697 => "00000000",
                     3698 => "01001010",
                     3699 => "00000101",
                     3700 => "00000000",
                     3701 => "01001010",
                     3702 => "01101000",
                     3703 => "00101010",
                     3704 => "10001000",
                     3705 => "11010000",
                     3706 => "11110001",
                     3707 => "10011101",
                     3708 => "11111100",
                     3709 => "00000110",
                     3710 => "01001000",
                     3711 => "00101001",
                     3712 => "00110000",
                     3713 => "00111101",
                     3714 => "01001010",
                     3715 => "00000111",
                     3716 => "11110000",
                     3717 => "00000111",
                     3718 => "01101000",
                     3719 => "00101001",
                     3720 => "11001111",
                     3721 => "10011101",
                     3722 => "11111100",
                     3723 => "00000110",
                     3724 => "01100000",
                     3725 => "01101000",
                     3726 => "10011101",
                     3727 => "01001010",
                     3728 => "00000111",
                     3729 => "01100000",
                     3730 => "10001101",
                     3731 => "00000110",
                     3732 => "00100000",
                     3733 => "11001000",
                     3734 => "10110001",
                     3735 => "00000000",
                     3736 => "10001101",
                     3737 => "00000110",
                     3738 => "00100000",
                     3739 => "11001000",
                     3740 => "10110001",
                     3741 => "00000000",
                     3742 => "00001010",
                     3743 => "01001000",
                     3744 => "10101101",
                     3745 => "01111000",
                     3746 => "00000111",
                     3747 => "00001001",
                     3748 => "00000100",
                     3749 => "10110000",
                     3750 => "00000010",
                     3751 => "00101001",
                     3752 => "11111011",
                     3753 => "00100000",
                     3754 => "11101101",
                     3755 => "10001110",
                     3756 => "01101000",
                     3757 => "00001010",
                     3758 => "10010000",
                     3759 => "00000011",
                     3760 => "00001001",
                     3761 => "00000010",
                     3762 => "11001000",
                     3763 => "01001010",
                     3764 => "01001010",
                     3765 => "10101010",
                     3766 => "10110000",
                     3767 => "00000001",
                     3768 => "11001000",
                     3769 => "10110001",
                     3770 => "00000000",
                     3771 => "10001101",
                     3772 => "00000111",
                     3773 => "00100000",
                     3774 => "11001010",
                     3775 => "11010000",
                     3776 => "11110101",
                     3777 => "00111000",
                     3778 => "10011000",
                     3779 => "01100101",
                     3780 => "00000000",
                     3781 => "10000101",
                     3782 => "00000000",
                     3783 => "10101001",
                     3784 => "00000000",
                     3785 => "01100101",
                     3786 => "00000001",
                     3787 => "10000101",
                     3788 => "00000001",
                     3789 => "10101001",
                     3790 => "00111111",
                     3791 => "10001101",
                     3792 => "00000110",
                     3793 => "00100000",
                     3794 => "10101001",
                     3795 => "00000000",
                     3796 => "10001101",
                     3797 => "00000110",
                     3798 => "00100000",
                     3799 => "10001101",
                     3800 => "00000110",
                     3801 => "00100000",
                     3802 => "10001101",
                     3803 => "00000110",
                     3804 => "00100000",
                     3805 => "10101110",
                     3806 => "00000010",
                     3807 => "00100000",
                     3808 => "10100000",
                     3809 => "00000000",
                     3810 => "10110001",
                     3811 => "00000000",
                     3812 => "11010000",
                     3813 => "10101100",
                     3814 => "10001101",
                     3815 => "00000101",
                     3816 => "00100000",
                     3817 => "10001101",
                     3818 => "00000101",
                     3819 => "00100000",
                     3820 => "01100000",
                     3821 => "10001101",
                     3822 => "00000000",
                     3823 => "00100000",
                     3824 => "10001101",
                     3825 => "01111000",
                     3826 => "00000111",
                     3827 => "01100000",
                     3828 => "11110000",
                     3829 => "00000110",
                     3830 => "01100010",
                     3831 => "00000110",
                     3832 => "01100010",
                     3833 => "00000110",
                     3834 => "01101101",
                     3835 => "00000010",
                     3836 => "01101101",
                     3837 => "00000010",
                     3838 => "01111010",
                     3839 => "00000011",
                     3840 => "00000110",
                     3841 => "00001100",
                     3842 => "00010010",
                     3843 => "00011000",
                     3844 => "00011110",
                     3845 => "00100100",
                     3846 => "10000101",
                     3847 => "00000000",
                     3848 => "00100000",
                     3849 => "00010001",
                     3850 => "10001111",
                     3851 => "10100101",
                     3852 => "00000000",
                     3853 => "01001010",
                     3854 => "01001010",
                     3855 => "01001010",
                     3856 => "01001010",
                     3857 => "00011000",
                     3858 => "01101001",
                     3859 => "00000001",
                     3860 => "00101001",
                     3861 => "00001111",
                     3862 => "11001001",
                     3863 => "00000110",
                     3864 => "10110000",
                     3865 => "01000100",
                     3866 => "01001000",
                     3867 => "00001010",
                     3868 => "10101000",
                     3869 => "10101110",
                     3870 => "00000000",
                     3871 => "00000011",
                     3872 => "10101001",
                     3873 => "00100000",
                     3874 => "11000000",
                     3875 => "00000000",
                     3876 => "11010000",
                     3877 => "00000010",
                     3878 => "10101001",
                     3879 => "00100010",
                     3880 => "10011101",
                     3881 => "00000001",
                     3882 => "00000011",
                     3883 => "10111001",
                     3884 => "11110100",
                     3885 => "10001110",
                     3886 => "10011101",
                     3887 => "00000010",
                     3888 => "00000011",
                     3889 => "10111001",
                     3890 => "11110101",
                     3891 => "10001110",
                     3892 => "10011101",
                     3893 => "00000011",
                     3894 => "00000011",
                     3895 => "10000101",
                     3896 => "00000011",
                     3897 => "10000110",
                     3898 => "00000010",
                     3899 => "01101000",
                     3900 => "10101010",
                     3901 => "10111101",
                     3902 => "00000000",
                     3903 => "10001111",
                     3904 => "00111000",
                     3905 => "11111001",
                     3906 => "11110101",
                     3907 => "10001110",
                     3908 => "10101000",
                     3909 => "10100110",
                     3910 => "00000010",
                     3911 => "10111001",
                     3912 => "11010111",
                     3913 => "00000111",
                     3914 => "10011101",
                     3915 => "00000100",
                     3916 => "00000011",
                     3917 => "11101000",
                     3918 => "11001000",
                     3919 => "11000110",
                     3920 => "00000011",
                     3921 => "11010000",
                     3922 => "11110100",
                     3923 => "10101001",
                     3924 => "00000000",
                     3925 => "10011101",
                     3926 => "00000100",
                     3927 => "00000011",
                     3928 => "11101000",
                     3929 => "11101000",
                     3930 => "11101000",
                     3931 => "10001110",
                     3932 => "00000000",
                     3933 => "00000011",
                     3934 => "01100000",
                     3935 => "10101101",
                     3936 => "01110000",
                     3937 => "00000111",
                     3938 => "11001001",
                     3939 => "00000000",
                     3940 => "11110000",
                     3941 => "00010110",
                     3942 => "10100010",
                     3943 => "00000101",
                     3944 => "10111101",
                     3945 => "00110100",
                     3946 => "00000001",
                     3947 => "00011000",
                     3948 => "01111001",
                     3949 => "11010111",
                     3950 => "00000111",
                     3951 => "00110000",
                     3952 => "00010110",
                     3953 => "11001001",
                     3954 => "00001010",
                     3955 => "10110000",
                     3956 => "00011001",
                     3957 => "10011001",
                     3958 => "11010111",
                     3959 => "00000111",
                     3960 => "10001000",
                     3961 => "11001010",
                     3962 => "00010000",
                     3963 => "11101100",
                     3964 => "10101001",
                     3965 => "00000000",
                     3966 => "10100010",
                     3967 => "00000110",
                     3968 => "10011101",
                     3969 => "00110011",
                     3970 => "00000001",
                     3971 => "11001010",
                     3972 => "00010000",
                     3973 => "11111010",
                     3974 => "01100000",
                     3975 => "11011110",
                     3976 => "00110011",
                     3977 => "00000001",
                     3978 => "10101001",
                     3979 => "00001001",
                     3980 => "11010000",
                     3981 => "11100111",
                     3982 => "00111000",
                     3983 => "11101001",
                     3984 => "00001010",
                     3985 => "11111110",
                     3986 => "00110011",
                     3987 => "00000001",
                     3988 => "01001100",
                     3989 => "01110101",
                     3990 => "10001111",
                     3991 => "10100010",
                     3992 => "00000101",
                     3993 => "00100000",
                     3994 => "10011110",
                     3995 => "10001111",
                     3996 => "10100010",
                     3997 => "00001011",
                     3998 => "10100000",
                     3999 => "00000101",
                     4000 => "00111000",
                     4001 => "10111101",
                     4002 => "11011101",
                     4003 => "00000111",
                     4004 => "11111001",
                     4005 => "11010111",
                     4006 => "00000111",
                     4007 => "11001010",
                     4008 => "10001000",
                     4009 => "00010000",
                     4010 => "11110110",
                     4011 => "10010000",
                     4012 => "00001110",
                     4013 => "11101000",
                     4014 => "11001000",
                     4015 => "10111101",
                     4016 => "11011101",
                     4017 => "00000111",
                     4018 => "10011001",
                     4019 => "11010111",
                     4020 => "00000111",
                     4021 => "11101000",
                     4022 => "11001000",
                     4023 => "11000000",
                     4024 => "00000110",
                     4025 => "10010000",
                     4026 => "11110100",
                     4027 => "01100000",
                     4028 => "00000100",
                     4029 => "00110000",
                     4030 => "01001000",
                     4031 => "01100000",
                     4032 => "01111000",
                     4033 => "10010000",
                     4034 => "10101000",
                     4035 => "11000000",
                     4036 => "11011000",
                     4037 => "11101000",
                     4038 => "00100100",
                     4039 => "11111000",
                     4040 => "11111100",
                     4041 => "00101000",
                     4042 => "00101100",
                     4043 => "00011000",
                     4044 => "11111111",
                     4045 => "00100011",
                     4046 => "01011000",
                     4047 => "10100000",
                     4048 => "01101111",
                     4049 => "00100000",
                     4050 => "11001100",
                     4051 => "10010000",
                     4052 => "10100000",
                     4053 => "00011111",
                     4054 => "10011001",
                     4055 => "10110000",
                     4056 => "00000111",
                     4057 => "10001000",
                     4058 => "00010000",
                     4059 => "11111010",
                     4060 => "10101001",
                     4061 => "00011000",
                     4062 => "10001101",
                     4063 => "10100010",
                     4064 => "00000111",
                     4065 => "00100000",
                     4066 => "00000011",
                     4067 => "10011100",
                     4068 => "10100000",
                     4069 => "01001011",
                     4070 => "00100000",
                     4071 => "11001100",
                     4072 => "10010000",
                     4073 => "10100010",
                     4074 => "00100001",
                     4075 => "10101001",
                     4076 => "00000000",
                     4077 => "10011101",
                     4078 => "10000000",
                     4079 => "00000111",
                     4080 => "11001010",
                     4081 => "00010000",
                     4082 => "11111010",
                     4083 => "10101101",
                     4084 => "01011011",
                     4085 => "00000111",
                     4086 => "10101100",
                     4087 => "01010010",
                     4088 => "00000111",
                     4089 => "11110000",
                     4090 => "00000011",
                     4091 => "10101101",
                     4092 => "01010001",
                     4093 => "00000111",
                     4094 => "10001101",
                     4095 => "00011010",
                     4096 => "00000111",
                     4097 => "10001101",
                     4098 => "00100101",
                     4099 => "00000111",
                     4100 => "10001101",
                     4101 => "00101000",
                     4102 => "00000111",
                     4103 => "00100000",
                     4104 => "00111000",
                     4105 => "10110000",
                     4106 => "10100000",
                     4107 => "00100000",
                     4108 => "00101001",
                     4109 => "00000001",
                     4110 => "11110000",
                     4111 => "00000010",
                     4112 => "10100000",
                     4113 => "00100100",
                     4114 => "10001100",
                     4115 => "00100000",
                     4116 => "00000111",
                     4117 => "10100000",
                     4118 => "10000000",
                     4119 => "10001100",
                     4120 => "00100001",
                     4121 => "00000111",
                     4122 => "00001010",
                     4123 => "00001010",
                     4124 => "00001010",
                     4125 => "00001010",
                     4126 => "10001101",
                     4127 => "10100000",
                     4128 => "00000110",
                     4129 => "11001110",
                     4130 => "00110000",
                     4131 => "00000111",
                     4132 => "11001110",
                     4133 => "00110001",
                     4134 => "00000111",
                     4135 => "11001110",
                     4136 => "00110010",
                     4137 => "00000111",
                     4138 => "10101001",
                     4139 => "00001011",
                     4140 => "10001101",
                     4141 => "00011110",
                     4142 => "00000111",
                     4143 => "00100000",
                     4144 => "00100010",
                     4145 => "10011100",
                     4146 => "10101101",
                     4147 => "01101010",
                     4148 => "00000111",
                     4149 => "11010000",
                     4150 => "00010000",
                     4151 => "10101101",
                     4152 => "01011111",
                     4153 => "00000111",
                     4154 => "11001001",
                     4155 => "00000100",
                     4156 => "10010000",
                     4157 => "00001100",
                     4158 => "11010000",
                     4159 => "00000111",
                     4160 => "10101101",
                     4161 => "01011100",
                     4162 => "00000111",
                     4163 => "11001001",
                     4164 => "00000010",
                     4165 => "10010000",
                     4166 => "00000011",
                     4167 => "11101110",
                     4168 => "11001100",
                     4169 => "00000110",
                     4170 => "10101101",
                     4171 => "01011011",
                     4172 => "00000111",
                     4173 => "11110000",
                     4174 => "00000101",
                     4175 => "10101001",
                     4176 => "00000010",
                     4177 => "10001101",
                     4178 => "00010000",
                     4179 => "00000111",
                     4180 => "10101001",
                     4181 => "10000000",
                     4182 => "10000101",
                     4183 => "11111011",
                     4184 => "10101001",
                     4185 => "00000001",
                     4186 => "10001101",
                     4187 => "01110100",
                     4188 => "00000111",
                     4189 => "11101110",
                     4190 => "01110010",
                     4191 => "00000111",
                     4192 => "01100000",
                     4193 => "10101001",
                     4194 => "00000001",
                     4195 => "10001101",
                     4196 => "01010111",
                     4197 => "00000111",
                     4198 => "10001101",
                     4199 => "01010100",
                     4200 => "00000111",
                     4201 => "10101001",
                     4202 => "00000010",
                     4203 => "10001101",
                     4204 => "01011010",
                     4205 => "00000111",
                     4206 => "10001101",
                     4207 => "01100001",
                     4208 => "00000111",
                     4209 => "10101001",
                     4210 => "00000000",
                     4211 => "10001101",
                     4212 => "01110100",
                     4213 => "00000111",
                     4214 => "10101000",
                     4215 => "10011001",
                     4216 => "00000000",
                     4217 => "00000011",
                     4218 => "11001000",
                     4219 => "11010000",
                     4220 => "11111010",
                     4221 => "10001101",
                     4222 => "01011001",
                     4223 => "00000111",
                     4224 => "10001101",
                     4225 => "01101001",
                     4226 => "00000111",
                     4227 => "10001101",
                     4228 => "00101000",
                     4229 => "00000111",
                     4230 => "10101001",
                     4231 => "11111111",
                     4232 => "10001101",
                     4233 => "10100000",
                     4234 => "00000011",
                     4235 => "10101101",
                     4236 => "00011010",
                     4237 => "00000111",
                     4238 => "01001110",
                     4239 => "01111000",
                     4240 => "00000111",
                     4241 => "00101001",
                     4242 => "00000001",
                     4243 => "01101010",
                     4244 => "00101110",
                     4245 => "01111000",
                     4246 => "00000111",
                     4247 => "00100000",
                     4248 => "11101101",
                     4249 => "10010000",
                     4250 => "10101001",
                     4251 => "00111000",
                     4252 => "10001101",
                     4253 => "11100011",
                     4254 => "00000110",
                     4255 => "10101001",
                     4256 => "01001000",
                     4257 => "10001101",
                     4258 => "11100010",
                     4259 => "00000110",
                     4260 => "10101001",
                     4261 => "01011000",
                     4262 => "10001101",
                     4263 => "11100001",
                     4264 => "00000110",
                     4265 => "10100010",
                     4266 => "00001110",
                     4267 => "10111101",
                     4268 => "10111100",
                     4269 => "10001111",
                     4270 => "10011101",
                     4271 => "11100100",
                     4272 => "00000110",
                     4273 => "11001010",
                     4274 => "00010000",
                     4275 => "11110111",
                     4276 => "10100000",
                     4277 => "00000011",
                     4278 => "10111001",
                     4279 => "11001011",
                     4280 => "10001111",
                     4281 => "10011001",
                     4282 => "00000000",
                     4283 => "00000010",
                     4284 => "10001000",
                     4285 => "00010000",
                     4286 => "11110111",
                     4287 => "00100000",
                     4288 => "10101111",
                     4289 => "10010010",
                     4290 => "00100000",
                     4291 => "10101010",
                     4292 => "10010010",
                     4293 => "11101110",
                     4294 => "00100010",
                     4295 => "00000111",
                     4296 => "11101110",
                     4297 => "01110010",
                     4298 => "00000111",
                     4299 => "01100000",
                     4300 => "10100010",
                     4301 => "00000111",
                     4302 => "10101001",
                     4303 => "00000000",
                     4304 => "10000101",
                     4305 => "00000110",
                     4306 => "10000110",
                     4307 => "00000111",
                     4308 => "11100000",
                     4309 => "00000001",
                     4310 => "11010000",
                     4311 => "00000100",
                     4312 => "11000000",
                     4313 => "01100000",
                     4314 => "10110000",
                     4315 => "00000010",
                     4316 => "10010001",
                     4317 => "00000110",
                     4318 => "10001000",
                     4319 => "11000000",
                     4320 => "11111111",
                     4321 => "11010000",
                     4322 => "11110001",
                     4323 => "11001010",
                     4324 => "00010000",
                     4325 => "11101100",
                     4326 => "01100000",
                     4327 => "00000010",
                     4328 => "00000001",
                     4329 => "00000100",
                     4330 => "00001000",
                     4331 => "00010000",
                     4332 => "00100000",
                     4333 => "10101101",
                     4334 => "01110000",
                     4335 => "00000111",
                     4336 => "11110000",
                     4337 => "00100011",
                     4338 => "10101101",
                     4339 => "01010010",
                     4340 => "00000111",
                     4341 => "11001001",
                     4342 => "00000010",
                     4343 => "11110000",
                     4344 => "00001101",
                     4345 => "10100000",
                     4346 => "00000101",
                     4347 => "10101101",
                     4348 => "00010000",
                     4349 => "00000111",
                     4350 => "11001001",
                     4351 => "00000110",
                     4352 => "11110000",
                     4353 => "00001110",
                     4354 => "11001001",
                     4355 => "00000111",
                     4356 => "11110000",
                     4357 => "00001010",
                     4358 => "10101100",
                     4359 => "01001110",
                     4360 => "00000111",
                     4361 => "10101101",
                     4362 => "01000011",
                     4363 => "00000111",
                     4364 => "11110000",
                     4365 => "00000010",
                     4366 => "10100000",
                     4367 => "00000100",
                     4368 => "10111001",
                     4369 => "11100111",
                     4370 => "10010000",
                     4371 => "10000101",
                     4372 => "11111011",
                     4373 => "01100000",
                     4374 => "00101000",
                     4375 => "00011000",
                     4376 => "00111000",
                     4377 => "00101000",
                     4378 => "00001000",
                     4379 => "00000000",
                     4380 => "00000000",
                     4381 => "00100000",
                     4382 => "10110000",
                     4383 => "01010000",
                     4384 => "00000000",
                     4385 => "00000000",
                     4386 => "10110000",
                     4387 => "10110000",
                     4388 => "11110000",
                     4389 => "00000000",
                     4390 => "00100000",
                     4391 => "00000000",
                     4392 => "00000000",
                     4393 => "00000000",
                     4394 => "00000000",
                     4395 => "00000000",
                     4396 => "00000000",
                     4397 => "00100000",
                     4398 => "00000100",
                     4399 => "00000011",
                     4400 => "00000010",
                     4401 => "10101101",
                     4402 => "00011010",
                     4403 => "00000111",
                     4404 => "10000101",
                     4405 => "01101101",
                     4406 => "10101001",
                     4407 => "01110000",
                     4408 => "10001101",
                     4409 => "00001010",
                     4410 => "00000111",
                     4411 => "10101001",
                     4412 => "00000001",
                     4413 => "10000101",
                     4414 => "00110011",
                     4415 => "10000101",
                     4416 => "10110101",
                     4417 => "10101001",
                     4418 => "00000000",
                     4419 => "10000101",
                     4420 => "00011101",
                     4421 => "11001110",
                     4422 => "10010000",
                     4423 => "00000100",
                     4424 => "10100000",
                     4425 => "00000000",
                     4426 => "10001100",
                     4427 => "01011011",
                     4428 => "00000111",
                     4429 => "10101101",
                     4430 => "01001110",
                     4431 => "00000111",
                     4432 => "11010000",
                     4433 => "00000001",
                     4434 => "11001000",
                     4435 => "10001100",
                     4436 => "00000100",
                     4437 => "00000111",
                     4438 => "10101110",
                     4439 => "00010000",
                     4440 => "00000111",
                     4441 => "10101100",
                     4442 => "01010010",
                     4443 => "00000111",
                     4444 => "11110000",
                     4445 => "00000111",
                     4446 => "11000000",
                     4447 => "00000001",
                     4448 => "11110000",
                     4449 => "00000011",
                     4450 => "10111110",
                     4451 => "00011000",
                     4452 => "10010001",
                     4453 => "10111001",
                     4454 => "00010110",
                     4455 => "10010001",
                     4456 => "10000101",
                     4457 => "10000110",
                     4458 => "10111101",
                     4459 => "00011100",
                     4460 => "10010001",
                     4461 => "10000101",
                     4462 => "11001110",
                     4463 => "10111101",
                     4464 => "00100101",
                     4465 => "10010001",
                     4466 => "10001101",
                     4467 => "11000100",
                     4468 => "00000011",
                     4469 => "00100000",
                     4470 => "11110001",
                     4471 => "10000101",
                     4472 => "10101100",
                     4473 => "00010101",
                     4474 => "00000111",
                     4475 => "11110000",
                     4476 => "00011010",
                     4477 => "10101101",
                     4478 => "01010111",
                     4479 => "00000111",
                     4480 => "11110000",
                     4481 => "00010101",
                     4482 => "10111001",
                     4483 => "00101101",
                     4484 => "10010001",
                     4485 => "10001101",
                     4486 => "11111000",
                     4487 => "00000111",
                     4488 => "10101001",
                     4489 => "00000001",
                     4490 => "10001101",
                     4491 => "11111010",
                     4492 => "00000111",
                     4493 => "01001010",
                     4494 => "10001101",
                     4495 => "11111001",
                     4496 => "00000111",
                     4497 => "10001101",
                     4498 => "01010111",
                     4499 => "00000111",
                     4500 => "10001101",
                     4501 => "10011111",
                     4502 => "00000111",
                     4503 => "10101100",
                     4504 => "01011000",
                     4505 => "00000111",
                     4506 => "11110000",
                     4507 => "00010100",
                     4508 => "10101001",
                     4509 => "00000011",
                     4510 => "10000101",
                     4511 => "00011101",
                     4512 => "10100010",
                     4513 => "00000000",
                     4514 => "00100000",
                     4515 => "10001001",
                     4516 => "10111101",
                     4517 => "10101001",
                     4518 => "11110000",
                     4519 => "10000101",
                     4520 => "11010111",
                     4521 => "10100010",
                     4522 => "00000101",
                     4523 => "10100000",
                     4524 => "00000000",
                     4525 => "00100000",
                     4526 => "00100011",
                     4527 => "10111001",
                     4528 => "10101100",
                     4529 => "01001110",
                     4530 => "00000111",
                     4531 => "11010000",
                     4532 => "00000011",
                     4533 => "00100000",
                     4534 => "00001011",
                     4535 => "10110111",
                     4536 => "10101001",
                     4537 => "00000111",
                     4538 => "10000101",
                     4539 => "00001110",
                     4540 => "01100000",
                     4541 => "01010110",
                     4542 => "01000000",
                     4543 => "01100101",
                     4544 => "01110000",
                     4545 => "01100110",
                     4546 => "01000000",
                     4547 => "01100110",
                     4548 => "01000000",
                     4549 => "01100110",
                     4550 => "01000000",
                     4551 => "01100110",
                     4552 => "01100000",
                     4553 => "01100101",
                     4554 => "01110000",
                     4555 => "00000000",
                     4556 => "00000000",
                     4557 => "11101110",
                     4558 => "01110100",
                     4559 => "00000111",
                     4560 => "10101001",
                     4561 => "00000000",
                     4562 => "10001101",
                     4563 => "00100010",
                     4564 => "00000111",
                     4565 => "10101001",
                     4566 => "10000000",
                     4567 => "10000101",
                     4568 => "11111100",
                     4569 => "11001110",
                     4570 => "01011010",
                     4571 => "00000111",
                     4572 => "00010000",
                     4573 => "00001011",
                     4574 => "10101001",
                     4575 => "00000000",
                     4576 => "10001101",
                     4577 => "01110010",
                     4578 => "00000111",
                     4579 => "10101001",
                     4580 => "00000011",
                     4581 => "10001101",
                     4582 => "01110000",
                     4583 => "00000111",
                     4584 => "01100000",
                     4585 => "10101101",
                     4586 => "01011111",
                     4587 => "00000111",
                     4588 => "00001010",
                     4589 => "10101010",
                     4590 => "10101101",
                     4591 => "01011100",
                     4592 => "00000111",
                     4593 => "00101001",
                     4594 => "00000010",
                     4595 => "11110000",
                     4596 => "00000001",
                     4597 => "11101000",
                     4598 => "10111100",
                     4599 => "10111101",
                     4600 => "10010001",
                     4601 => "10101101",
                     4602 => "01011100",
                     4603 => "00000111",
                     4604 => "01001010",
                     4605 => "10011000",
                     4606 => "10110000",
                     4607 => "00000100",
                     4608 => "01001010",
                     4609 => "01001010",
                     4610 => "01001010",
                     4611 => "01001010",
                     4612 => "00101001",
                     4613 => "00001111",
                     4614 => "11001101",
                     4615 => "00011010",
                     4616 => "00000111",
                     4617 => "11110000",
                     4618 => "00000100",
                     4619 => "10010000",
                     4620 => "00000010",
                     4621 => "10101001",
                     4622 => "00000000",
                     4623 => "10001101",
                     4624 => "01011011",
                     4625 => "00000111",
                     4626 => "00100000",
                     4627 => "10000010",
                     4628 => "10010010",
                     4629 => "01001100",
                     4630 => "01100100",
                     4631 => "10010010",
                     4632 => "10101101",
                     4633 => "01110010",
                     4634 => "00000111",
                     4635 => "00100000",
                     4636 => "00000100",
                     4637 => "10001110",
                     4638 => "00100100",
                     4639 => "10010010",
                     4640 => "01100111",
                     4641 => "10000101",
                     4642 => "00110111",
                     4643 => "10010010",
                     4644 => "10101001",
                     4645 => "00000000",
                     4646 => "10001101",
                     4647 => "00111100",
                     4648 => "00000111",
                     4649 => "10001101",
                     4650 => "00100010",
                     4651 => "00000111",
                     4652 => "10101001",
                     4653 => "00000010",
                     4654 => "10000101",
                     4655 => "11111100",
                     4656 => "11101110",
                     4657 => "01110100",
                     4658 => "00000111",
                     4659 => "11101110",
                     4660 => "01110010",
                     4661 => "00000111",
                     4662 => "01100000",
                     4663 => "10101001",
                     4664 => "00000000",
                     4665 => "10001101",
                     4666 => "01110100",
                     4667 => "00000111",
                     4668 => "10101101",
                     4669 => "11111100",
                     4670 => "00000110",
                     4671 => "00101001",
                     4672 => "00010000",
                     4673 => "11010000",
                     4674 => "00000101",
                     4675 => "10101101",
                     4676 => "10100000",
                     4677 => "00000111",
                     4678 => "11010000",
                     4679 => "00111001",
                     4680 => "10101001",
                     4681 => "10000000",
                     4682 => "10000101",
                     4683 => "11111100",
                     4684 => "00100000",
                     4685 => "10000010",
                     4686 => "10010010",
                     4687 => "10010000",
                     4688 => "00010011",
                     4689 => "10101101",
                     4690 => "01011111",
                     4691 => "00000111",
                     4692 => "10001101",
                     4693 => "11111101",
                     4694 => "00000111",
                     4695 => "10101001",
                     4696 => "00000000",
                     4697 => "00001010",
                     4698 => "10001101",
                     4699 => "01110010",
                     4700 => "00000111",
                     4701 => "10001101",
                     4702 => "10100000",
                     4703 => "00000111",
                     4704 => "10001101",
                     4705 => "01110000",
                     4706 => "00000111",
                     4707 => "01100000",
                     4708 => "00100000",
                     4709 => "00000011",
                     4710 => "10011100",
                     4711 => "10101001",
                     4712 => "00000001",
                     4713 => "10001101",
                     4714 => "01010100",
                     4715 => "00000111",
                     4716 => "11101110",
                     4717 => "01010111",
                     4718 => "00000111",
                     4719 => "10101001",
                     4720 => "00000000",
                     4721 => "10001101",
                     4722 => "01000111",
                     4723 => "00000111",
                     4724 => "10001101",
                     4725 => "01010110",
                     4726 => "00000111",
                     4727 => "10000101",
                     4728 => "00001110",
                     4729 => "10001101",
                     4730 => "01110010",
                     4731 => "00000111",
                     4732 => "10101001",
                     4733 => "00000001",
                     4734 => "10001101",
                     4735 => "01110000",
                     4736 => "00000111",
                     4737 => "01100000",
                     4738 => "00111000",
                     4739 => "10101101",
                     4740 => "01111010",
                     4741 => "00000111",
                     4742 => "11110000",
                     4743 => "00100001",
                     4744 => "10101101",
                     4745 => "01100001",
                     4746 => "00000111",
                     4747 => "00110000",
                     4748 => "00011100",
                     4749 => "10101101",
                     4750 => "01010011",
                     4751 => "00000111",
                     4752 => "01001001",
                     4753 => "00000001",
                     4754 => "10001101",
                     4755 => "01010011",
                     4756 => "00000111",
                     4757 => "10100010",
                     4758 => "00000110",
                     4759 => "10111101",
                     4760 => "01011010",
                     4761 => "00000111",
                     4762 => "01001000",
                     4763 => "10111101",
                     4764 => "01100001",
                     4765 => "00000111",
                     4766 => "10011101",
                     4767 => "01011010",
                     4768 => "00000111",
                     4769 => "01101000",
                     4770 => "10011101",
                     4771 => "01100001",
                     4772 => "00000111",
                     4773 => "11001010",
                     4774 => "00010000",
                     4775 => "11101111",
                     4776 => "00011000",
                     4777 => "01100000",
                     4778 => "10101001",
                     4779 => "11111111",
                     4780 => "10001101",
                     4781 => "11001001",
                     4782 => "00000110",
                     4783 => "01100000",
                     4784 => "10101100",
                     4785 => "00011111",
                     4786 => "00000111",
                     4787 => "11010000",
                     4788 => "00000101",
                     4789 => "10100000",
                     4790 => "00001000",
                     4791 => "10001100",
                     4792 => "00011111",
                     4793 => "00000111",
                     4794 => "10001000",
                     4795 => "10011000",
                     4796 => "00100000",
                     4797 => "11001000",
                     4798 => "10010010",
                     4799 => "11001110",
                     4800 => "00011111",
                     4801 => "00000111",
                     4802 => "11010000",
                     4803 => "00000011",
                     4804 => "00100000",
                     4805 => "01101010",
                     4806 => "10001001",
                     4807 => "01100000",
                     4808 => "00100000",
                     4809 => "00000100",
                     4810 => "10001110",
                     4811 => "11011011",
                     4812 => "10010010",
                     4813 => "10101110",
                     4814 => "10001000",
                     4815 => "10101110",
                     4816 => "10001000",
                     4817 => "11111100",
                     4818 => "10010011",
                     4819 => "11011011",
                     4820 => "10010010",
                     4821 => "10101110",
                     4822 => "10001000",
                     4823 => "10101110",
                     4824 => "10001000",
                     4825 => "11111100",
                     4826 => "10010011",
                     4827 => "11101110",
                     4828 => "00100110",
                     4829 => "00000111",
                     4830 => "10101101",
                     4831 => "00100110",
                     4832 => "00000111",
                     4833 => "00101001",
                     4834 => "00001111",
                     4835 => "11010000",
                     4836 => "00000110",
                     4837 => "10001101",
                     4838 => "00100110",
                     4839 => "00000111",
                     4840 => "11101110",
                     4841 => "00100101",
                     4842 => "00000111",
                     4843 => "11101110",
                     4844 => "10100000",
                     4845 => "00000110",
                     4846 => "10101101",
                     4847 => "10100000",
                     4848 => "00000110",
                     4849 => "00101001",
                     4850 => "00011111",
                     4851 => "10001101",
                     4852 => "10100000",
                     4853 => "00000110",
                     4854 => "01100000",
                     4855 => "00000000",
                     4856 => "00110000",
                     4857 => "01100000",
                     4858 => "10010011",
                     4859 => "00000000",
                     4860 => "00000000",
                     4861 => "00010001",
                     4862 => "00010010",
                     4863 => "00010010",
                     4864 => "00010011",
                     4865 => "00000000",
                     4866 => "00000000",
                     4867 => "01010001",
                     4868 => "01010010",
                     4869 => "01010011",
                     4870 => "00000000",
                     4871 => "00000000",
                     4872 => "00000000",
                     4873 => "00000000",
                     4874 => "00000000",
                     4875 => "00000000",
                     4876 => "00000001",
                     4877 => "00000010",
                     4878 => "00000010",
                     4879 => "00000011",
                     4880 => "00000000",
                     4881 => "00000000",
                     4882 => "00000000",
                     4883 => "00000000",
                     4884 => "00000000",
                     4885 => "00000000",
                     4886 => "10010001",
                     4887 => "10010010",
                     4888 => "10010011",
                     4889 => "00000000",
                     4890 => "00000000",
                     4891 => "00000000",
                     4892 => "00000000",
                     4893 => "01010001",
                     4894 => "01010010",
                     4895 => "01010011",
                     4896 => "01000001",
                     4897 => "01000010",
                     4898 => "01000011",
                     4899 => "00000000",
                     4900 => "00000000",
                     4901 => "00000000",
                     4902 => "00000000",
                     4903 => "00000000",
                     4904 => "10010001",
                     4905 => "10010010",
                     4906 => "10010111",
                     4907 => "10000111",
                     4908 => "10001000",
                     4909 => "10001001",
                     4910 => "10011001",
                     4911 => "00000000",
                     4912 => "00000000",
                     4913 => "00000000",
                     4914 => "00010001",
                     4915 => "00010010",
                     4916 => "00010011",
                     4917 => "10100100",
                     4918 => "10100101",
                     4919 => "10100101",
                     4920 => "10100101",
                     4921 => "10100110",
                     4922 => "10010111",
                     4923 => "10011000",
                     4924 => "10011001",
                     4925 => "00000001",
                     4926 => "00000010",
                     4927 => "00000011",
                     4928 => "00000000",
                     4929 => "10100100",
                     4930 => "10100101",
                     4931 => "10100110",
                     4932 => "00000000",
                     4933 => "00010001",
                     4934 => "00010010",
                     4935 => "00010010",
                     4936 => "00010010",
                     4937 => "00010011",
                     4938 => "00000000",
                     4939 => "00000000",
                     4940 => "00000000",
                     4941 => "00000000",
                     4942 => "00000001",
                     4943 => "00000010",
                     4944 => "00000010",
                     4945 => "00000011",
                     4946 => "00000000",
                     4947 => "10100100",
                     4948 => "10100101",
                     4949 => "10100101",
                     4950 => "10100110",
                     4951 => "00000000",
                     4952 => "00000000",
                     4953 => "00000000",
                     4954 => "00010001",
                     4955 => "00010010",
                     4956 => "00010010",
                     4957 => "00010011",
                     4958 => "00000000",
                     4959 => "00000000",
                     4960 => "00000000",
                     4961 => "00000000",
                     4962 => "00000000",
                     4963 => "00000000",
                     4964 => "00000000",
                     4965 => "10011100",
                     4966 => "00000000",
                     4967 => "10001011",
                     4968 => "10101010",
                     4969 => "10101010",
                     4970 => "10101010",
                     4971 => "10101010",
                     4972 => "00010001",
                     4973 => "00010010",
                     4974 => "00010011",
                     4975 => "10001011",
                     4976 => "00000000",
                     4977 => "10011100",
                     4978 => "10011100",
                     4979 => "00000000",
                     4980 => "00000000",
                     4981 => "00000001",
                     4982 => "00000010",
                     4983 => "00000011",
                     4984 => "00010001",
                     4985 => "00010010",
                     4986 => "00010010",
                     4987 => "00010011",
                     4988 => "00000000",
                     4989 => "00000000",
                     4990 => "00000000",
                     4991 => "00000000",
                     4992 => "10101010",
                     4993 => "10101010",
                     4994 => "10011100",
                     4995 => "10101010",
                     4996 => "00000000",
                     4997 => "10001011",
                     4998 => "00000000",
                     4999 => "00000001",
                     5000 => "00000010",
                     5001 => "00000011",
                     5002 => "10000000",
                     5003 => "10000011",
                     5004 => "00000000",
                     5005 => "10000001",
                     5006 => "10000100",
                     5007 => "00000000",
                     5008 => "10000010",
                     5009 => "10000101",
                     5010 => "00000000",
                     5011 => "00000010",
                     5012 => "00000000",
                     5013 => "00000000",
                     5014 => "00000011",
                     5015 => "00000000",
                     5016 => "00000000",
                     5017 => "00000100",
                     5018 => "00000000",
                     5019 => "00000000",
                     5020 => "00000000",
                     5021 => "00000101",
                     5022 => "00000110",
                     5023 => "00000111",
                     5024 => "00000110",
                     5025 => "00001010",
                     5026 => "00000000",
                     5027 => "00001000",
                     5028 => "00001001",
                     5029 => "01001101",
                     5030 => "00000000",
                     5031 => "00000000",
                     5032 => "00001101",
                     5033 => "00001111",
                     5034 => "01001110",
                     5035 => "00001110",
                     5036 => "01001110",
                     5037 => "01001110",
                     5038 => "00000000",
                     5039 => "00001101",
                     5040 => "00011010",
                     5041 => "10000110",
                     5042 => "10000111",
                     5043 => "10000111",
                     5044 => "10000111",
                     5045 => "10000111",
                     5046 => "10000111",
                     5047 => "10000111",
                     5048 => "10000111",
                     5049 => "10000111",
                     5050 => "10000111",
                     5051 => "10000111",
                     5052 => "01101001",
                     5053 => "01101001",
                     5054 => "00000000",
                     5055 => "00000000",
                     5056 => "00000000",
                     5057 => "00000000",
                     5058 => "00000000",
                     5059 => "01000101",
                     5060 => "01000111",
                     5061 => "01000111",
                     5062 => "01000111",
                     5063 => "01000111",
                     5064 => "01000111",
                     5065 => "00000000",
                     5066 => "00000000",
                     5067 => "00000000",
                     5068 => "00000000",
                     5069 => "00000000",
                     5070 => "00000000",
                     5071 => "00000000",
                     5072 => "00000000",
                     5073 => "00000000",
                     5074 => "00000000",
                     5075 => "00000000",
                     5076 => "00000000",
                     5077 => "00000000",
                     5078 => "10000110",
                     5079 => "10000111",
                     5080 => "01101001",
                     5081 => "01010100",
                     5082 => "01010010",
                     5083 => "01100010",
                     5084 => "00000000",
                     5085 => "00000000",
                     5086 => "00000000",
                     5087 => "00011000",
                     5088 => "00000001",
                     5089 => "00011000",
                     5090 => "00000111",
                     5091 => "00011000",
                     5092 => "00001111",
                     5093 => "00011000",
                     5094 => "11111111",
                     5095 => "00011000",
                     5096 => "00000001",
                     5097 => "00011111",
                     5098 => "00000111",
                     5099 => "00011111",
                     5100 => "00001111",
                     5101 => "00011111",
                     5102 => "10000001",
                     5103 => "00011111",
                     5104 => "00000001",
                     5105 => "00000000",
                     5106 => "10001111",
                     5107 => "00011111",
                     5108 => "11110001",
                     5109 => "00011111",
                     5110 => "11111001",
                     5111 => "00011000",
                     5112 => "11110001",
                     5113 => "00011000",
                     5114 => "11111111",
                     5115 => "00011111",
                     5116 => "10101101",
                     5117 => "00101000",
                     5118 => "00000111",
                     5119 => "11110000",
                     5120 => "00000011",
                     5121 => "00100000",
                     5122 => "00001000",
                     5123 => "10010101",
                     5124 => "10100010",
                     5125 => "00001100",
                     5126 => "10101001",
                     5127 => "00000000",
                     5128 => "10011101",
                     5129 => "10100001",
                     5130 => "00000110",
                     5131 => "11001010",
                     5132 => "00010000",
                     5133 => "11111010",
                     5134 => "10101100",
                     5135 => "01000010",
                     5136 => "00000111",
                     5137 => "11110000",
                     5138 => "01000010",
                     5139 => "10101101",
                     5140 => "00100101",
                     5141 => "00000111",
                     5142 => "11001001",
                     5143 => "00000011",
                     5144 => "00110000",
                     5145 => "00000101",
                     5146 => "00111000",
                     5147 => "11101001",
                     5148 => "00000011",
                     5149 => "00010000",
                     5150 => "11110111",
                     5151 => "00001010",
                     5152 => "00001010",
                     5153 => "00001010",
                     5154 => "00001010",
                     5155 => "01111001",
                     5156 => "11110110",
                     5157 => "10010010",
                     5158 => "01101101",
                     5159 => "00100110",
                     5160 => "00000111",
                     5161 => "10101010",
                     5162 => "10111101",
                     5163 => "11111010",
                     5164 => "10010010",
                     5165 => "11110000",
                     5166 => "00100110",
                     5167 => "01001000",
                     5168 => "00101001",
                     5169 => "00001111",
                     5170 => "00111000",
                     5171 => "11101001",
                     5172 => "00000001",
                     5173 => "10000101",
                     5174 => "00000000",
                     5175 => "00001010",
                     5176 => "01100101",
                     5177 => "00000000",
                     5178 => "10101010",
                     5179 => "01101000",
                     5180 => "01001010",
                     5181 => "01001010",
                     5182 => "01001010",
                     5183 => "01001010",
                     5184 => "10101000",
                     5185 => "10101001",
                     5186 => "00000011",
                     5187 => "10000101",
                     5188 => "00000000",
                     5189 => "10111101",
                     5190 => "10001010",
                     5191 => "10010011",
                     5192 => "10011001",
                     5193 => "10100001",
                     5194 => "00000110",
                     5195 => "11101000",
                     5196 => "11001000",
                     5197 => "11000000",
                     5198 => "00001011",
                     5199 => "11110000",
                     5200 => "00000100",
                     5201 => "11000110",
                     5202 => "00000000",
                     5203 => "11010000",
                     5204 => "11110000",
                     5205 => "10101110",
                     5206 => "01000001",
                     5207 => "00000111",
                     5208 => "11110000",
                     5209 => "00010011",
                     5210 => "10111100",
                     5211 => "10101101",
                     5212 => "10010011",
                     5213 => "10100010",
                     5214 => "00000000",
                     5215 => "10111001",
                     5216 => "10110001",
                     5217 => "10010011",
                     5218 => "11110000",
                     5219 => "00000011",
                     5220 => "10011101",
                     5221 => "10100001",
                     5222 => "00000110",
                     5223 => "11001000",
                     5224 => "11101000",
                     5225 => "11100000",
                     5226 => "00001101",
                     5227 => "11010000",
                     5228 => "11110010",
                     5229 => "10101100",
                     5230 => "01001110",
                     5231 => "00000111",
                     5232 => "11010000",
                     5233 => "00001100",
                     5234 => "10101101",
                     5235 => "01011111",
                     5236 => "00000111",
                     5237 => "11001001",
                     5238 => "00000111",
                     5239 => "11010000",
                     5240 => "00000101",
                     5241 => "10101001",
                     5242 => "01100010",
                     5243 => "01001100",
                     5244 => "10001000",
                     5245 => "10010100",
                     5246 => "10111001",
                     5247 => "11011000",
                     5248 => "10010011",
                     5249 => "10101100",
                     5250 => "01000011",
                     5251 => "00000111",
                     5252 => "11110000",
                     5253 => "00000010",
                     5254 => "10101001",
                     5255 => "10001000",
                     5256 => "10000101",
                     5257 => "00000111",
                     5258 => "10100010",
                     5259 => "00000000",
                     5260 => "10101101",
                     5261 => "00100111",
                     5262 => "00000111",
                     5263 => "00001010",
                     5264 => "10101000",
                     5265 => "10111001",
                     5266 => "11011100",
                     5267 => "10010011",
                     5268 => "10000101",
                     5269 => "00000000",
                     5270 => "11001000",
                     5271 => "10000100",
                     5272 => "00000001",
                     5273 => "10101101",
                     5274 => "01000011",
                     5275 => "00000111",
                     5276 => "11110000",
                     5277 => "00001010",
                     5278 => "11100000",
                     5279 => "00000000",
                     5280 => "11110000",
                     5281 => "00000110",
                     5282 => "10100101",
                     5283 => "00000000",
                     5284 => "00101001",
                     5285 => "00001000",
                     5286 => "10000101",
                     5287 => "00000000",
                     5288 => "10100000",
                     5289 => "00000000",
                     5290 => "10111001",
                     5291 => "10010000",
                     5292 => "11000110",
                     5293 => "00100100",
                     5294 => "00000000",
                     5295 => "11110000",
                     5296 => "00000101",
                     5297 => "10100101",
                     5298 => "00000111",
                     5299 => "10011101",
                     5300 => "10100001",
                     5301 => "00000110",
                     5302 => "11101000",
                     5303 => "11100000",
                     5304 => "00001101",
                     5305 => "11110000",
                     5306 => "00011000",
                     5307 => "10101101",
                     5308 => "01001110",
                     5309 => "00000111",
                     5310 => "11001001",
                     5311 => "00000010",
                     5312 => "11010000",
                     5313 => "00001000",
                     5314 => "11100000",
                     5315 => "00001011",
                     5316 => "11010000",
                     5317 => "00000100",
                     5318 => "10101001",
                     5319 => "01010100",
                     5320 => "10000101",
                     5321 => "00000111",
                     5322 => "11001000",
                     5323 => "11000000",
                     5324 => "00001000",
                     5325 => "11010000",
                     5326 => "11011011",
                     5327 => "10100100",
                     5328 => "00000001",
                     5329 => "11010000",
                     5330 => "10111110",
                     5331 => "00100000",
                     5332 => "00001000",
                     5333 => "10010101",
                     5334 => "10101101",
                     5335 => "10100000",
                     5336 => "00000110",
                     5337 => "00100000",
                     5338 => "11100011",
                     5339 => "10011011",
                     5340 => "10100010",
                     5341 => "00000000",
                     5342 => "10100000",
                     5343 => "00000000",
                     5344 => "10000100",
                     5345 => "00000000",
                     5346 => "10111101",
                     5347 => "10100001",
                     5348 => "00000110",
                     5349 => "00101001",
                     5350 => "11000000",
                     5351 => "00001010",
                     5352 => "00101010",
                     5353 => "00101010",
                     5354 => "10101000",
                     5355 => "10111101",
                     5356 => "10100001",
                     5357 => "00000110",
                     5358 => "11011001",
                     5359 => "00000100",
                     5360 => "10010101",
                     5361 => "10110000",
                     5362 => "00000010",
                     5363 => "10101001",
                     5364 => "00000000",
                     5365 => "10100100",
                     5366 => "00000000",
                     5367 => "10010001",
                     5368 => "00000110",
                     5369 => "10011000",
                     5370 => "00011000",
                     5371 => "01101001",
                     5372 => "00010000",
                     5373 => "10101000",
                     5374 => "11101000",
                     5375 => "11100000",
                     5376 => "00001101",
                     5377 => "10010000",
                     5378 => "11011101",
                     5379 => "01100000",
                     5380 => "00010000",
                     5381 => "01010001",
                     5382 => "10001000",
                     5383 => "11000000",
                     5384 => "10100010",
                     5385 => "00000010",
                     5386 => "10000110",
                     5387 => "00001000",
                     5388 => "10101001",
                     5389 => "00000000",
                     5390 => "10001101",
                     5391 => "00101001",
                     5392 => "00000111",
                     5393 => "10101100",
                     5394 => "00101100",
                     5395 => "00000111",
                     5396 => "10110001",
                     5397 => "11100111",
                     5398 => "11001001",
                     5399 => "11111101",
                     5400 => "11110000",
                     5401 => "01001011",
                     5402 => "10111101",
                     5403 => "00110000",
                     5404 => "00000111",
                     5405 => "00010000",
                     5406 => "01000110",
                     5407 => "11001000",
                     5408 => "10110001",
                     5409 => "11100111",
                     5410 => "00001010",
                     5411 => "10010000",
                     5412 => "00001011",
                     5413 => "10101101",
                     5414 => "00101011",
                     5415 => "00000111",
                     5416 => "11010000",
                     5417 => "00000110",
                     5418 => "11101110",
                     5419 => "00101011",
                     5420 => "00000111",
                     5421 => "11101110",
                     5422 => "00101010",
                     5423 => "00000111",
                     5424 => "10001000",
                     5425 => "10110001",
                     5426 => "11100111",
                     5427 => "00101001",
                     5428 => "00001111",
                     5429 => "11001001",
                     5430 => "00001101",
                     5431 => "11010000",
                     5432 => "00011011",
                     5433 => "11001000",
                     5434 => "10110001",
                     5435 => "11100111",
                     5436 => "10001000",
                     5437 => "00101001",
                     5438 => "01000000",
                     5439 => "11010000",
                     5440 => "00011100",
                     5441 => "10101101",
                     5442 => "00101011",
                     5443 => "00000111",
                     5444 => "11010000",
                     5445 => "00010111",
                     5446 => "11001000",
                     5447 => "10110001",
                     5448 => "11100111",
                     5449 => "00101001",
                     5450 => "00011111",
                     5451 => "10001101",
                     5452 => "00101010",
                     5453 => "00000111",
                     5454 => "11101110",
                     5455 => "00101011",
                     5456 => "00000111",
                     5457 => "01001100",
                     5458 => "01101110",
                     5459 => "10010101",
                     5460 => "11001001",
                     5461 => "00001110",
                     5462 => "11010000",
                     5463 => "00000101",
                     5464 => "10101101",
                     5465 => "00101000",
                     5466 => "00000111",
                     5467 => "11010000",
                     5468 => "00001000",
                     5469 => "10101101",
                     5470 => "00101010",
                     5471 => "00000111",
                     5472 => "11001101",
                     5473 => "00100101",
                     5474 => "00000111",
                     5475 => "10010000",
                     5476 => "00000110",
                     5477 => "00100000",
                     5478 => "10010101",
                     5479 => "10010101",
                     5480 => "01001100",
                     5481 => "01110001",
                     5482 => "10010101",
                     5483 => "11101110",
                     5484 => "00101001",
                     5485 => "00000111",
                     5486 => "00100000",
                     5487 => "10001001",
                     5488 => "10010101",
                     5489 => "10100110",
                     5490 => "00001000",
                     5491 => "10111101",
                     5492 => "00110000",
                     5493 => "00000111",
                     5494 => "00110000",
                     5495 => "00000011",
                     5496 => "11011110",
                     5497 => "00110000",
                     5498 => "00000111",
                     5499 => "11001010",
                     5500 => "00010000",
                     5501 => "10001100",
                     5502 => "10101101",
                     5503 => "00101001",
                     5504 => "00000111",
                     5505 => "11010000",
                     5506 => "10000101",
                     5507 => "10101101",
                     5508 => "00101000",
                     5509 => "00000111",
                     5510 => "11010000",
                     5511 => "10000000",
                     5512 => "01100000",
                     5513 => "11101110",
                     5514 => "00101100",
                     5515 => "00000111",
                     5516 => "11101110",
                     5517 => "00101100",
                     5518 => "00000111",
                     5519 => "10101001",
                     5520 => "00000000",
                     5521 => "10001101",
                     5522 => "00101011",
                     5523 => "00000111",
                     5524 => "01100000",
                     5525 => "10111101",
                     5526 => "00110000",
                     5527 => "00000111",
                     5528 => "00110000",
                     5529 => "00000011",
                     5530 => "10111100",
                     5531 => "00101101",
                     5532 => "00000111",
                     5533 => "10100010",
                     5534 => "00010000",
                     5535 => "10110001",
                     5536 => "11100111",
                     5537 => "11001001",
                     5538 => "11111101",
                     5539 => "11110000",
                     5540 => "11100011",
                     5541 => "00101001",
                     5542 => "00001111",
                     5543 => "11001001",
                     5544 => "00001111",
                     5545 => "11110000",
                     5546 => "00001000",
                     5547 => "10100010",
                     5548 => "00001000",
                     5549 => "11001001",
                     5550 => "00001100",
                     5551 => "11110000",
                     5552 => "00000010",
                     5553 => "10100010",
                     5554 => "00000000",
                     5555 => "10000110",
                     5556 => "00000111",
                     5557 => "10100110",
                     5558 => "00001000",
                     5559 => "11001001",
                     5560 => "00001110",
                     5561 => "11010000",
                     5562 => "00001000",
                     5563 => "10101001",
                     5564 => "00000000",
                     5565 => "10000101",
                     5566 => "00000111",
                     5567 => "10101001",
                     5568 => "00101110",
                     5569 => "11010000",
                     5570 => "01010011",
                     5571 => "11001001",
                     5572 => "00001101",
                     5573 => "11010000",
                     5574 => "00011011",
                     5575 => "10101001",
                     5576 => "00100010",
                     5577 => "10000101",
                     5578 => "00000111",
                     5579 => "11001000",
                     5580 => "10110001",
                     5581 => "11100111",
                     5582 => "00101001",
                     5583 => "01000000",
                     5584 => "11110000",
                     5585 => "01100011",
                     5586 => "10110001",
                     5587 => "11100111",
                     5588 => "00101001",
                     5589 => "01111111",
                     5590 => "11001001",
                     5591 => "01001011",
                     5592 => "11010000",
                     5593 => "00000011",
                     5594 => "11101110",
                     5595 => "01000101",
                     5596 => "00000111",
                     5597 => "00101001",
                     5598 => "00111111",
                     5599 => "01001100",
                     5600 => "00010110",
                     5601 => "10010110",
                     5602 => "11001001",
                     5603 => "00001100",
                     5604 => "10110000",
                     5605 => "00100111",
                     5606 => "11001000",
                     5607 => "10110001",
                     5608 => "11100111",
                     5609 => "00101001",
                     5610 => "01110000",
                     5611 => "11010000",
                     5612 => "00001011",
                     5613 => "10101001",
                     5614 => "00010110",
                     5615 => "10000101",
                     5616 => "00000111",
                     5617 => "10110001",
                     5618 => "11100111",
                     5619 => "00101001",
                     5620 => "00001111",
                     5621 => "01001100",
                     5622 => "00010110",
                     5623 => "10010110",
                     5624 => "10000101",
                     5625 => "00000000",
                     5626 => "11001001",
                     5627 => "01110000",
                     5628 => "11010000",
                     5629 => "00001010",
                     5630 => "10110001",
                     5631 => "11100111",
                     5632 => "00101001",
                     5633 => "00001000",
                     5634 => "11110000",
                     5635 => "00000100",
                     5636 => "10101001",
                     5637 => "00000000",
                     5638 => "10000101",
                     5639 => "00000000",
                     5640 => "10100101",
                     5641 => "00000000",
                     5642 => "01001100",
                     5643 => "00010010",
                     5644 => "10010110",
                     5645 => "11001000",
                     5646 => "10110001",
                     5647 => "11100111",
                     5648 => "00101001",
                     5649 => "01110000",
                     5650 => "01001010",
                     5651 => "01001010",
                     5652 => "01001010",
                     5653 => "01001010",
                     5654 => "10000101",
                     5655 => "00000000",
                     5656 => "10111101",
                     5657 => "00110000",
                     5658 => "00000111",
                     5659 => "00010000",
                     5660 => "01000010",
                     5661 => "10101101",
                     5662 => "00101010",
                     5663 => "00000111",
                     5664 => "11001101",
                     5665 => "00100101",
                     5666 => "00000111",
                     5667 => "11110000",
                     5668 => "00010001",
                     5669 => "10101100",
                     5670 => "00101100",
                     5671 => "00000111",
                     5672 => "10110001",
                     5673 => "11100111",
                     5674 => "00101001",
                     5675 => "00001111",
                     5676 => "11001001",
                     5677 => "00001110",
                     5678 => "11010000",
                     5679 => "00000101",
                     5680 => "10101101",
                     5681 => "00101000",
                     5682 => "00000111",
                     5683 => "11010000",
                     5684 => "00100001",
                     5685 => "01100000",
                     5686 => "10101101",
                     5687 => "00101000",
                     5688 => "00000111",
                     5689 => "11110000",
                     5690 => "00001011",
                     5691 => "10101001",
                     5692 => "00000000",
                     5693 => "10001101",
                     5694 => "00101000",
                     5695 => "00000111",
                     5696 => "10001101",
                     5697 => "00101001",
                     5698 => "00000111",
                     5699 => "10000101",
                     5700 => "00001000",
                     5701 => "01100000",
                     5702 => "10101100",
                     5703 => "00101100",
                     5704 => "00000111",
                     5705 => "10110001",
                     5706 => "11100111",
                     5707 => "00101001",
                     5708 => "11110000",
                     5709 => "01001010",
                     5710 => "01001010",
                     5711 => "01001010",
                     5712 => "01001010",
                     5713 => "11001101",
                     5714 => "00100110",
                     5715 => "00000111",
                     5716 => "11010000",
                     5717 => "11011111",
                     5718 => "10101101",
                     5719 => "00101100",
                     5720 => "00000111",
                     5721 => "10011101",
                     5722 => "00101101",
                     5723 => "00000111",
                     5724 => "00100000",
                     5725 => "10001001",
                     5726 => "10010101",
                     5727 => "10100101",
                     5728 => "00000000",
                     5729 => "00011000",
                     5730 => "01100101",
                     5731 => "00000111",
                     5732 => "00100000",
                     5733 => "00000100",
                     5734 => "10001110",
                     5735 => "11100101",
                     5736 => "10011000",
                     5737 => "01000000",
                     5738 => "10010111",
                     5739 => "00101110",
                     5740 => "10011010",
                     5741 => "00111110",
                     5742 => "10011010",
                     5743 => "11110010",
                     5744 => "10011001",
                     5745 => "01010000",
                     5746 => "10011010",
                     5747 => "01011001",
                     5748 => "10011010",
                     5749 => "11100101",
                     5750 => "10011000",
                     5751 => "01000011",
                     5752 => "10011011",
                     5753 => "10111010",
                     5754 => "10010111",
                     5755 => "01111001",
                     5756 => "10011001",
                     5757 => "01111100",
                     5758 => "10011001",
                     5759 => "01111111",
                     5760 => "10011001",
                     5761 => "01010111",
                     5762 => "10011001",
                     5763 => "01101000",
                     5764 => "10011001",
                     5765 => "01101011",
                     5766 => "10011001",
                     5767 => "11010000",
                     5768 => "10011001",
                     5769 => "11010111",
                     5770 => "10011001",
                     5771 => "00000110",
                     5772 => "10011000",
                     5773 => "10110111",
                     5774 => "10011010",
                     5775 => "10101011",
                     5776 => "10011000",
                     5777 => "10010100",
                     5778 => "10011001",
                     5779 => "00010000",
                     5780 => "10011011",
                     5781 => "00010000",
                     5782 => "10011011",
                     5783 => "00010000",
                     5784 => "10011011",
                     5785 => "00000011",
                     5786 => "10011011",
                     5787 => "00011011",
                     5788 => "10011011",
                     5789 => "00011011",
                     5790 => "10011011",
                     5791 => "00011011",
                     5792 => "10011011",
                     5793 => "00010110",
                     5794 => "10011011",
                     5795 => "00011011",
                     5796 => "10011011",
                     5797 => "01101111",
                     5798 => "10011000",
                     5799 => "00011001",
                     5800 => "10011010",
                     5801 => "11010011",
                     5802 => "10011010",
                     5803 => "10000010",
                     5804 => "10011000",
                     5805 => "10011110",
                     5806 => "10011001",
                     5807 => "00001001",
                     5808 => "10011010",
                     5809 => "00001110",
                     5810 => "10011010",
                     5811 => "00000001",
                     5812 => "10011010",
                     5813 => "11110010",
                     5814 => "10010110",
                     5815 => "00001101",
                     5816 => "10010111",
                     5817 => "00001101",
                     5818 => "10010111",
                     5819 => "00101011",
                     5820 => "10010111",
                     5821 => "00101011",
                     5822 => "10010111",
                     5823 => "00101011",
                     5824 => "10010111",
                     5825 => "01000101",
                     5826 => "10010110",
                     5827 => "11000101",
                     5828 => "10010110",
                     5829 => "10111100",
                     5830 => "00101101",
                     5831 => "00000111",
                     5832 => "11001000",
                     5833 => "10110001",
                     5834 => "11100111",
                     5835 => "01001000",
                     5836 => "00101001",
                     5837 => "01000000",
                     5838 => "11010000",
                     5839 => "00010010",
                     5840 => "01101000",
                     5841 => "01001000",
                     5842 => "00101001",
                     5843 => "00001111",
                     5844 => "10001101",
                     5845 => "00100111",
                     5846 => "00000111",
                     5847 => "01101000",
                     5848 => "00101001",
                     5849 => "00110000",
                     5850 => "01001010",
                     5851 => "01001010",
                     5852 => "01001010",
                     5853 => "01001010",
                     5854 => "10001101",
                     5855 => "01000010",
                     5856 => "00000111",
                     5857 => "01100000",
                     5858 => "01101000",
                     5859 => "00101001",
                     5860 => "00000111",
                     5861 => "11001001",
                     5862 => "00000100",
                     5863 => "10010000",
                     5864 => "00000101",
                     5865 => "10001101",
                     5866 => "01000100",
                     5867 => "00000111",
                     5868 => "10101001",
                     5869 => "00000000",
                     5870 => "10001101",
                     5871 => "01000001",
                     5872 => "00000111",
                     5873 => "01100000",
                     5874 => "10100010",
                     5875 => "00000100",
                     5876 => "10101101",
                     5877 => "01011111",
                     5878 => "00000111",
                     5879 => "11110000",
                     5880 => "00001000",
                     5881 => "11101000",
                     5882 => "10101100",
                     5883 => "01001110",
                     5884 => "00000111",
                     5885 => "10001000",
                     5886 => "11010000",
                     5887 => "00000001",
                     5888 => "11101000",
                     5889 => "10001010",
                     5890 => "10001101",
                     5891 => "11010110",
                     5892 => "00000110",
                     5893 => "00100000",
                     5894 => "00001000",
                     5895 => "10001000",
                     5896 => "10101001",
                     5897 => "00001101",
                     5898 => "00100000",
                     5899 => "00010110",
                     5900 => "10010111",
                     5901 => "10101101",
                     5902 => "00100011",
                     5903 => "00000111",
                     5904 => "01001001",
                     5905 => "00000001",
                     5906 => "10001101",
                     5907 => "00100011",
                     5908 => "00000111",
                     5909 => "01100000",
                     5910 => "10000101",
                     5911 => "00000000",
                     5912 => "10101001",
                     5913 => "00000000",
                     5914 => "10100010",
                     5915 => "00000100",
                     5916 => "10110100",
                     5917 => "00010110",
                     5918 => "11000100",
                     5919 => "00000000",
                     5920 => "11010000",
                     5921 => "00000010",
                     5922 => "10010101",
                     5923 => "00001111",
                     5924 => "11001010",
                     5925 => "00010000",
                     5926 => "11110101",
                     5927 => "01100000",
                     5928 => "00010100",
                     5929 => "00010111",
                     5930 => "00011000",
                     5931 => "10100110",
                     5932 => "00000000",
                     5933 => "10111101",
                     5934 => "00100000",
                     5935 => "10010111",
                     5936 => "10100000",
                     5937 => "00000101",
                     5938 => "10001000",
                     5939 => "00110000",
                     5940 => "00000111",
                     5941 => "11011001",
                     5942 => "00010110",
                     5943 => "00000000",
                     5944 => "11010000",
                     5945 => "11111000",
                     5946 => "10101001",
                     5947 => "00000000",
                     5948 => "10001101",
                     5949 => "11001101",
                     5950 => "00000110",
                     5951 => "01100000",
                     5952 => "10101101",
                     5953 => "00110011",
                     5954 => "00000111",
                     5955 => "00100000",
                     5956 => "00000100",
                     5957 => "10001110",
                     5958 => "01001100",
                     5959 => "10010111",
                     5960 => "01111000",
                     5961 => "10010111",
                     5962 => "01101001",
                     5963 => "10011010",
                     5964 => "00100000",
                     5965 => "10111101",
                     5966 => "10011011",
                     5967 => "10111101",
                     5968 => "00110000",
                     5969 => "00000111",
                     5970 => "11110000",
                     5971 => "00011111",
                     5972 => "00010000",
                     5973 => "00010001",
                     5974 => "10011000",
                     5975 => "10011101",
                     5976 => "00110000",
                     5977 => "00000111",
                     5978 => "10101101",
                     5979 => "00100101",
                     5980 => "00000111",
                     5981 => "00001101",
                     5982 => "00100110",
                     5983 => "00000111",
                     5984 => "11110000",
                     5985 => "00000101",
                     5986 => "10101001",
                     5987 => "00010110",
                     5988 => "01001100",
                     5989 => "10110000",
                     5990 => "10010111",
                     5991 => "10100110",
                     5992 => "00000111",
                     5993 => "10101001",
                     5994 => "00010111",
                     5995 => "10011101",
                     5996 => "10100001",
                     5997 => "00000110",
                     5998 => "10101001",
                     5999 => "01001100",
                     6000 => "01001100",
                     6001 => "10101010",
                     6002 => "10010111",
                     6003 => "10101001",
                     6004 => "00011000",
                     6005 => "01001100",
                     6006 => "10110000",
                     6007 => "10010111",
                     6008 => "00100000",
                     6009 => "10101110",
                     6010 => "10011011",
                     6011 => "10000100",
                     6012 => "00000110",
                     6013 => "10010000",
                     6014 => "00001100",
                     6015 => "10111101",
                     6016 => "00110000",
                     6017 => "00000111",
                     6018 => "01001010",
                     6019 => "10011101",
                     6020 => "00110110",
                     6021 => "00000111",
                     6022 => "10101001",
                     6023 => "00011001",
                     6024 => "01001100",
                     6025 => "10110000",
                     6026 => "10010111",
                     6027 => "10101001",
                     6028 => "00011011",
                     6029 => "10111100",
                     6030 => "00110000",
                     6031 => "00000111",
                     6032 => "11110000",
                     6033 => "00011110",
                     6034 => "10111101",
                     6035 => "00110110",
                     6036 => "00000111",
                     6037 => "10000101",
                     6038 => "00000110",
                     6039 => "10100110",
                     6040 => "00000111",
                     6041 => "10101001",
                     6042 => "00011010",
                     6043 => "10011101",
                     6044 => "10100001",
                     6045 => "00000110",
                     6046 => "11000100",
                     6047 => "00000110",
                     6048 => "11010000",
                     6049 => "00101100",
                     6050 => "11101000",
                     6051 => "10101001",
                     6052 => "01001111",
                     6053 => "10011101",
                     6054 => "10100001",
                     6055 => "00000110",
                     6056 => "10101001",
                     6057 => "01010000",
                     6058 => "11101000",
                     6059 => "10100000",
                     6060 => "00001111",
                     6061 => "01001100",
                     6062 => "01111111",
                     6063 => "10011011",
                     6064 => "10100110",
                     6065 => "00000111",
                     6066 => "10100000",
                     6067 => "00000000",
                     6068 => "01001100",
                     6069 => "01111111",
                     6070 => "10011011",
                     6071 => "01000010",
                     6072 => "01000001",
                     6073 => "01000011",
                     6074 => "00100000",
                     6075 => "10101110",
                     6076 => "10011011",
                     6077 => "10100000",
                     6078 => "00000000",
                     6079 => "10110000",
                     6080 => "00000111",
                     6081 => "11001000",
                     6082 => "10111101",
                     6083 => "00110000",
                     6084 => "00000111",
                     6085 => "11010000",
                     6086 => "00000001",
                     6087 => "11001000",
                     6088 => "10111001",
                     6089 => "10110111",
                     6090 => "10010111",
                     6091 => "10001101",
                     6092 => "10100001",
                     6093 => "00000110",
                     6094 => "01100000",
                     6095 => "00000000",
                     6096 => "01000101",
                     6097 => "01000101",
                     6098 => "01000101",
                     6099 => "00000000",
                     6100 => "00000000",
                     6101 => "01001000",
                     6102 => "01000111",
                     6103 => "01000110",
                     6104 => "00000000",
                     6105 => "01000101",
                     6106 => "01001001",
                     6107 => "01001001",
                     6108 => "01001001",
                     6109 => "01000101",
                     6110 => "01000111",
                     6111 => "01000111",
                     6112 => "01001010",
                     6113 => "01000111",
                     6114 => "01000111",
                     6115 => "01000111",
                     6116 => "01000111",
                     6117 => "01001011",
                     6118 => "01000111",
                     6119 => "01000111",
                     6120 => "01001001",
                     6121 => "01001001",
                     6122 => "01001001",
                     6123 => "01001001",
                     6124 => "01001001",
                     6125 => "01000111",
                     6126 => "01001010",
                     6127 => "01000111",
                     6128 => "01001010",
                     6129 => "01000111",
                     6130 => "01000111",
                     6131 => "01001011",
                     6132 => "01000111",
                     6133 => "01001011",
                     6134 => "01000111",
                     6135 => "01000111",
                     6136 => "01000111",
                     6137 => "01000111",
                     6138 => "01000111",
                     6139 => "01000111",
                     6140 => "01001010",
                     6141 => "01000111",
                     6142 => "01001010",
                     6143 => "01000111",
                     6144 => "01001010",
                     6145 => "01001011",
                     6146 => "01000111",
                     6147 => "01001011",
                     6148 => "01000111",
                     6149 => "01001011",
                     6150 => "00100000",
                     6151 => "10111101",
                     6152 => "10011011",
                     6153 => "10000100",
                     6154 => "00000111",
                     6155 => "10100000",
                     6156 => "00000100",
                     6157 => "00100000",
                     6158 => "10110001",
                     6159 => "10011011",
                     6160 => "10001010",
                     6161 => "01001000",
                     6162 => "10111100",
                     6163 => "00110000",
                     6164 => "00000111",
                     6165 => "10100110",
                     6166 => "00000111",
                     6167 => "10101001",
                     6168 => "00001011",
                     6169 => "10000101",
                     6170 => "00000110",
                     6171 => "10111001",
                     6172 => "11001111",
                     6173 => "10010111",
                     6174 => "10011101",
                     6175 => "10100001",
                     6176 => "00000110",
                     6177 => "11101000",
                     6178 => "10100101",
                     6179 => "00000110",
                     6180 => "11110000",
                     6181 => "00000111",
                     6182 => "11001000",
                     6183 => "11001000",
                     6184 => "11001000",
                     6185 => "11001000",
                     6186 => "11001000",
                     6187 => "11000110",
                     6188 => "00000110",
                     6189 => "11100000",
                     6190 => "00001011",
                     6191 => "11010000",
                     6192 => "11101010",
                     6193 => "01101000",
                     6194 => "10101010",
                     6195 => "10101101",
                     6196 => "00100101",
                     6197 => "00000111",
                     6198 => "11110000",
                     6199 => "00110110",
                     6200 => "10111101",
                     6201 => "00110000",
                     6202 => "00000111",
                     6203 => "11001001",
                     6204 => "00000001",
                     6205 => "11110000",
                     6206 => "00101010",
                     6207 => "10100100",
                     6208 => "00000111",
                     6209 => "11010000",
                     6210 => "00000100",
                     6211 => "11001001",
                     6212 => "00000011",
                     6213 => "11110000",
                     6214 => "00100010",
                     6215 => "11001001",
                     6216 => "00000010",
                     6217 => "11010000",
                     6218 => "00100011",
                     6219 => "00100000",
                     6220 => "11001101",
                     6221 => "10011011",
                     6222 => "01001000",
                     6223 => "00100000",
                     6224 => "01001010",
                     6225 => "10011001",
                     6226 => "01101000",
                     6227 => "10010101",
                     6228 => "10000111",
                     6229 => "10101101",
                     6230 => "00100101",
                     6231 => "00000111",
                     6232 => "10010101",
                     6233 => "01101110",
                     6234 => "10101001",
                     6235 => "00000001",
                     6236 => "10010101",
                     6237 => "10110110",
                     6238 => "10010101",
                     6239 => "00001111",
                     6240 => "10101001",
                     6241 => "10010000",
                     6242 => "10010101",
                     6243 => "11001111",
                     6244 => "10101001",
                     6245 => "00110001",
                     6246 => "10010101",
                     6247 => "00010110",
                     6248 => "01100000",
                     6249 => "10100000",
                     6250 => "01010010",
                     6251 => "10001100",
                     6252 => "10101011",
                     6253 => "00000110",
                     6254 => "01100000",
                     6255 => "00100000",
                     6256 => "10111101",
                     6257 => "10011011",
                     6258 => "10111100",
                     6259 => "00110000",
                     6260 => "00000111",
                     6261 => "10100110",
                     6262 => "00000111",
                     6263 => "10101001",
                     6264 => "01101011",
                     6265 => "10011101",
                     6266 => "10100001",
                     6267 => "00000110",
                     6268 => "10101001",
                     6269 => "01101100",
                     6270 => "10011101",
                     6271 => "10100010",
                     6272 => "00000110",
                     6273 => "01100000",
                     6274 => "10100000",
                     6275 => "00000011",
                     6276 => "00100000",
                     6277 => "10110001",
                     6278 => "10011011",
                     6279 => "10100000",
                     6280 => "00001010",
                     6281 => "00100000",
                     6282 => "10110011",
                     6283 => "10011000",
                     6284 => "10110000",
                     6285 => "00010000",
                     6286 => "10100010",
                     6287 => "00000110",
                     6288 => "10101001",
                     6289 => "00000000",
                     6290 => "10011101",
                     6291 => "10100001",
                     6292 => "00000110",
                     6293 => "11001010",
                     6294 => "00010000",
                     6295 => "11111000",
                     6296 => "10111001",
                     6297 => "11011101",
                     6298 => "10011000",
                     6299 => "10001101",
                     6300 => "10101000",
                     6301 => "00000110",
                     6302 => "01100000",
                     6303 => "00010101",
                     6304 => "00010100",
                     6305 => "00000000",
                     6306 => "00000000",
                     6307 => "00010101",
                     6308 => "00011110",
                     6309 => "00011101",
                     6310 => "00011100",
                     6311 => "00010101",
                     6312 => "00100001",
                     6313 => "00100000",
                     6314 => "00011111",
                     6315 => "10100000",
                     6316 => "00000011",
                     6317 => "00100000",
                     6318 => "10110001",
                     6319 => "10011011",
                     6320 => "00100000",
                     6321 => "10111101",
                     6322 => "10011011",
                     6323 => "10001000",
                     6324 => "10001000",
                     6325 => "10000100",
                     6326 => "00000101",
                     6327 => "10111100",
                     6328 => "00110000",
                     6329 => "00000111",
                     6330 => "10000100",
                     6331 => "00000110",
                     6332 => "10100110",
                     6333 => "00000101",
                     6334 => "11101000",
                     6335 => "10111001",
                     6336 => "10011111",
                     6337 => "10011000",
                     6338 => "11001001",
                     6339 => "00000000",
                     6340 => "11110000",
                     6341 => "00001000",
                     6342 => "10100010",
                     6343 => "00000000",
                     6344 => "10100100",
                     6345 => "00000101",
                     6346 => "00100000",
                     6347 => "01111111",
                     6348 => "10011011",
                     6349 => "00011000",
                     6350 => "10100100",
                     6351 => "00000110",
                     6352 => "10111001",
                     6353 => "10100011",
                     6354 => "10011000",
                     6355 => "10011101",
                     6356 => "10100001",
                     6357 => "00000110",
                     6358 => "10111001",
                     6359 => "10100111",
                     6360 => "10011000",
                     6361 => "10011101",
                     6362 => "10100010",
                     6363 => "00000110",
                     6364 => "01100000",
                     6365 => "00010001",
                     6366 => "00010000",
                     6367 => "00010101",
                     6368 => "00010100",
                     6369 => "00010011",
                     6370 => "00010010",
                     6371 => "00010101",
                     6372 => "00010100",
                     6373 => "00100000",
                     6374 => "00111001",
                     6375 => "10011001",
                     6376 => "10100101",
                     6377 => "00000000",
                     6378 => "11110000",
                     6379 => "00000100",
                     6380 => "11001000",
                     6381 => "11001000",
                     6382 => "11001000",
                     6383 => "11001000",
                     6384 => "10011000",
                     6385 => "01001000",
                     6386 => "10101101",
                     6387 => "01100000",
                     6388 => "00000111",
                     6389 => "00001101",
                     6390 => "01011111",
                     6391 => "00000111",
                     6392 => "11110000",
                     6393 => "00101011",
                     6394 => "10111100",
                     6395 => "00110000",
                     6396 => "00000111",
                     6397 => "11110000",
                     6398 => "00100110",
                     6399 => "00100000",
                     6400 => "01001010",
                     6401 => "10011001",
                     6402 => "10110000",
                     6403 => "00100001",
                     6404 => "00100000",
                     6405 => "11001101",
                     6406 => "10011011",
                     6407 => "00011000",
                     6408 => "01101001",
                     6409 => "00001000",
                     6410 => "10010101",
                     6411 => "10000111",
                     6412 => "10101101",
                     6413 => "00100101",
                     6414 => "00000111",
                     6415 => "01101001",
                     6416 => "00000000",
                     6417 => "10010101",
                     6418 => "01101110",
                     6419 => "10101001",
                     6420 => "00000001",
                     6421 => "10010101",
                     6422 => "10110110",
                     6423 => "10010101",
                     6424 => "00001111",
                     6425 => "00100000",
                     6426 => "11010101",
                     6427 => "10011011",
                     6428 => "10010101",
                     6429 => "11001111",
                     6430 => "10101001",
                     6431 => "00001101",
                     6432 => "10010101",
                     6433 => "00010110",
                     6434 => "00100000",
                     6435 => "10001101",
                     6436 => "11000111",
                     6437 => "01101000",
                     6438 => "10101000",
                     6439 => "10100110",
                     6440 => "00000111",
                     6441 => "10111001",
                     6442 => "11011101",
                     6443 => "10011000",
                     6444 => "10011101",
                     6445 => "10100001",
                     6446 => "00000110",
                     6447 => "11101000",
                     6448 => "10111001",
                     6449 => "11011111",
                     6450 => "10011000",
                     6451 => "10100100",
                     6452 => "00000110",
                     6453 => "10001000",
                     6454 => "01001100",
                     6455 => "01111111",
                     6456 => "10011011",
                     6457 => "10100000",
                     6458 => "00000001",
                     6459 => "00100000",
                     6460 => "10110001",
                     6461 => "10011011",
                     6462 => "00100000",
                     6463 => "10111101",
                     6464 => "10011011",
                     6465 => "10011000",
                     6466 => "00101001",
                     6467 => "00000111",
                     6468 => "10000101",
                     6469 => "00000110",
                     6470 => "10111100",
                     6471 => "00110000",
                     6472 => "00000111",
                     6473 => "01100000",
                     6474 => "10100010",
                     6475 => "00000000",
                     6476 => "00011000",
                     6477 => "10110101",
                     6478 => "00001111",
                     6479 => "11110000",
                     6480 => "00000101",
                     6481 => "11101000",
                     6482 => "11100000",
                     6483 => "00000101",
                     6484 => "11010000",
                     6485 => "11110110",
                     6486 => "01100000",
                     6487 => "00100000",
                     6488 => "10101110",
                     6489 => "10011011",
                     6490 => "10101001",
                     6491 => "10000110",
                     6492 => "10001101",
                     6493 => "10101011",
                     6494 => "00000110",
                     6495 => "10100010",
                     6496 => "00001011",
                     6497 => "10100000",
                     6498 => "00000001",
                     6499 => "10101001",
                     6500 => "10000111",
                     6501 => "01001100",
                     6502 => "01111111",
                     6503 => "10011011",
                     6504 => "10101001",
                     6505 => "00000011",
                     6506 => "00101100",
                     6507 => "10101001",
                     6508 => "00000111",
                     6509 => "01001000",
                     6510 => "00100000",
                     6511 => "10101110",
                     6512 => "10011011",
                     6513 => "01101000",
                     6514 => "10101010",
                     6515 => "10101001",
                     6516 => "11000000",
                     6517 => "10011101",
                     6518 => "10100001",
                     6519 => "00000110",
                     6520 => "01100000",
                     6521 => "10101001",
                     6522 => "00000110",
                     6523 => "00101100",
                     6524 => "10101001",
                     6525 => "00000111",
                     6526 => "00101100",
                     6527 => "10101001",
                     6528 => "00001001",
                     6529 => "01001000",
                     6530 => "00100000",
                     6531 => "10101110",
                     6532 => "10011011",
                     6533 => "01101000",
                     6534 => "10101010",
                     6535 => "10101001",
                     6536 => "00001011",
                     6537 => "10011101",
                     6538 => "10100001",
                     6539 => "00000110",
                     6540 => "11101000",
                     6541 => "10100000",
                     6542 => "00000000",
                     6543 => "10101001",
                     6544 => "01100011",
                     6545 => "01001100",
                     6546 => "01111111",
                     6547 => "10011011",
                     6548 => "00100000",
                     6549 => "10111101",
                     6550 => "10011011",
                     6551 => "10100010",
                     6552 => "00000010",
                     6553 => "10101001",
                     6554 => "01101101",
                     6555 => "01001100",
                     6556 => "01111111",
                     6557 => "10011011",
                     6558 => "10101001",
                     6559 => "00100100",
                     6560 => "10001101",
                     6561 => "10100001",
                     6562 => "00000110",
                     6563 => "10100010",
                     6564 => "00000001",
                     6565 => "10100000",
                     6566 => "00001000",
                     6567 => "10101001",
                     6568 => "00100101",
                     6569 => "00100000",
                     6570 => "01111111",
                     6571 => "10011011",
                     6572 => "10101001",
                     6573 => "01100001",
                     6574 => "10001101",
                     6575 => "10101011",
                     6576 => "00000110",
                     6577 => "00100000",
                     6578 => "11001101",
                     6579 => "10011011",
                     6580 => "00111000",
                     6581 => "11101001",
                     6582 => "00001000",
                     6583 => "10000101",
                     6584 => "10001100",
                     6585 => "10101101",
                     6586 => "00100101",
                     6587 => "00000111",
                     6588 => "11101001",
                     6589 => "00000000",
                     6590 => "10000101",
                     6591 => "01110011",
                     6592 => "10101001",
                     6593 => "00110000",
                     6594 => "10000101",
                     6595 => "11010100",
                     6596 => "10101001",
                     6597 => "10110000",
                     6598 => "10001101",
                     6599 => "00001101",
                     6600 => "00000001",
                     6601 => "10101001",
                     6602 => "00110000",
                     6603 => "10000101",
                     6604 => "00011011",
                     6605 => "11100110",
                     6606 => "00010100",
                     6607 => "01100000",
                     6608 => "10100010",
                     6609 => "00000000",
                     6610 => "10100000",
                     6611 => "00001111",
                     6612 => "01001100",
                     6613 => "11101001",
                     6614 => "10011001",
                     6615 => "10001010",
                     6616 => "01001000",
                     6617 => "10100010",
                     6618 => "00000001",
                     6619 => "10100000",
                     6620 => "00001111",
                     6621 => "10101001",
                     6622 => "01000100",
                     6623 => "00100000",
                     6624 => "01111111",
                     6625 => "10011011",
                     6626 => "01101000",
                     6627 => "10101010",
                     6628 => "00100000",
                     6629 => "10111101",
                     6630 => "10011011",
                     6631 => "10100010",
                     6632 => "00000001",
                     6633 => "10101001",
                     6634 => "01000000",
                     6635 => "01001100",
                     6636 => "01111111",
                     6637 => "10011011",
                     6638 => "11000011",
                     6639 => "11000010",
                     6640 => "11000010",
                     6641 => "11000010",
                     6642 => "10101100",
                     6643 => "01001110",
                     6644 => "00000111",
                     6645 => "10111001",
                     6646 => "11101110",
                     6647 => "10011001",
                     6648 => "01001100",
                     6649 => "01000100",
                     6650 => "10011010",
                     6651 => "00000110",
                     6652 => "00000111",
                     6653 => "00001000",
                     6654 => "11000101",
                     6655 => "00001100",
                     6656 => "10001001",
                     6657 => "10100000",
                     6658 => "00001100",
                     6659 => "00100000",
                     6660 => "10110001",
                     6661 => "10011011",
                     6662 => "01001100",
                     6663 => "00001110",
                     6664 => "10011010",
                     6665 => "10101001",
                     6666 => "00001000",
                     6667 => "10001101",
                     6668 => "01110011",
                     6669 => "00000111",
                     6670 => "10100100",
                     6671 => "00000000",
                     6672 => "10111110",
                     6673 => "11111001",
                     6674 => "10011001",
                     6675 => "10111001",
                     6676 => "11111100",
                     6677 => "10011001",
                     6678 => "01001100",
                     6679 => "00100000",
                     6680 => "10011010",
                     6681 => "00100000",
                     6682 => "10111101",
                     6683 => "10011011",
                     6684 => "10100110",
                     6685 => "00000111",
                     6686 => "10101001",
                     6687 => "11000100",
                     6688 => "10100000",
                     6689 => "00000000",
                     6690 => "01001100",
                     6691 => "01111111",
                     6692 => "10011011",
                     6693 => "01101001",
                     6694 => "01100001",
                     6695 => "01100001",
                     6696 => "01100010",
                     6697 => "00100010",
                     6698 => "01010001",
                     6699 => "01010010",
                     6700 => "01010010",
                     6701 => "10001000",
                     6702 => "10101100",
                     6703 => "01001110",
                     6704 => "00000111",
                     6705 => "10101101",
                     6706 => "01000011",
                     6707 => "00000111",
                     6708 => "11110000",
                     6709 => "00000010",
                     6710 => "10100000",
                     6711 => "00000100",
                     6712 => "10111001",
                     6713 => "00101001",
                     6714 => "10011010",
                     6715 => "01001100",
                     6716 => "01000100",
                     6717 => "10011010",
                     6718 => "10101100",
                     6719 => "01001110",
                     6720 => "00000111",
                     6721 => "10111001",
                     6722 => "00100101",
                     6723 => "10011010",
                     6724 => "01001000",
                     6725 => "00100000",
                     6726 => "10101110",
                     6727 => "10011011",
                     6728 => "10100110",
                     6729 => "00000111",
                     6730 => "10100000",
                     6731 => "00000000",
                     6732 => "01101000",
                     6733 => "01001100",
                     6734 => "01111111",
                     6735 => "10011011",
                     6736 => "10101100",
                     6737 => "01001110",
                     6738 => "00000111",
                     6739 => "10111001",
                     6740 => "00101001",
                     6741 => "10011010",
                     6742 => "01001100",
                     6743 => "01011111",
                     6744 => "10011010",
                     6745 => "10101100",
                     6746 => "01001110",
                     6747 => "00000111",
                     6748 => "10111001",
                     6749 => "00100101",
                     6750 => "10011010",
                     6751 => "01001000",
                     6752 => "00100000",
                     6753 => "10111101",
                     6754 => "10011011",
                     6755 => "01101000",
                     6756 => "10100110",
                     6757 => "00000111",
                     6758 => "01001100",
                     6759 => "01111111",
                     6760 => "10011011",
                     6761 => "00100000",
                     6762 => "10111101",
                     6763 => "10011011",
                     6764 => "10100110",
                     6765 => "00000111",
                     6766 => "10101001",
                     6767 => "01100100",
                     6768 => "10011101",
                     6769 => "10100001",
                     6770 => "00000110",
                     6771 => "11101000",
                     6772 => "10001000",
                     6773 => "00110000",
                     6774 => "00001110",
                     6775 => "10101001",
                     6776 => "01100101",
                     6777 => "10011101",
                     6778 => "10100001",
                     6779 => "00000110",
                     6780 => "11101000",
                     6781 => "10001000",
                     6782 => "00110000",
                     6783 => "00000101",
                     6784 => "10101001",
                     6785 => "01100110",
                     6786 => "00100000",
                     6787 => "01111111",
                     6788 => "10011011",
                     6789 => "10101110",
                     6790 => "01101010",
                     6791 => "00000100",
                     6792 => "00100000",
                     6793 => "11010101",
                     6794 => "10011011",
                     6795 => "10011101",
                     6796 => "01110111",
                     6797 => "00000100",
                     6798 => "10101101",
                     6799 => "00100101",
                     6800 => "00000111",
                     6801 => "10011101",
                     6802 => "01101011",
                     6803 => "00000100",
                     6804 => "00100000",
                     6805 => "11001101",
                     6806 => "10011011",
                     6807 => "10011101",
                     6808 => "01110001",
                     6809 => "00000100",
                     6810 => "11101000",
                     6811 => "11100000",
                     6812 => "00000110",
                     6813 => "10010000",
                     6814 => "00000010",
                     6815 => "10100010",
                     6816 => "00000000",
                     6817 => "10001110",
                     6818 => "01101010",
                     6819 => "00000100",
                     6820 => "01100000",
                     6821 => "00000111",
                     6822 => "00000111",
                     6823 => "00000110",
                     6824 => "00000101",
                     6825 => "00000100",
                     6826 => "00000011",
                     6827 => "00000010",
                     6828 => "00000001",
                     6829 => "00000000",
                     6830 => "00000011",
                     6831 => "00000011",
                     6832 => "00000100",
                     6833 => "00000101",
                     6834 => "00000110",
                     6835 => "00000111",
                     6836 => "00001000",
                     6837 => "00001001",
                     6838 => "00001010",
                     6839 => "00100000",
                     6840 => "10101110",
                     6841 => "10011011",
                     6842 => "10010000",
                     6843 => "00000101",
                     6844 => "10101001",
                     6845 => "00001001",
                     6846 => "10001101",
                     6847 => "00110100",
                     6848 => "00000111",
                     6849 => "11001110",
                     6850 => "00110100",
                     6851 => "00000111",
                     6852 => "10101100",
                     6853 => "00110100",
                     6854 => "00000111",
                     6855 => "10111110",
                     6856 => "10101110",
                     6857 => "10011010",
                     6858 => "10111001",
                     6859 => "10100101",
                     6860 => "10011010",
                     6861 => "10101000",
                     6862 => "10101001",
                     6863 => "01100001",
                     6864 => "01001100",
                     6865 => "01111111",
                     6866 => "10011011",
                     6867 => "00100000",
                     6868 => "10111101",
                     6869 => "10011011",
                     6870 => "00100000",
                     6871 => "01001010",
                     6872 => "10011001",
                     6873 => "10110000",
                     6874 => "00100111",
                     6875 => "00100000",
                     6876 => "11001101",
                     6877 => "10011011",
                     6878 => "10010101",
                     6879 => "10000111",
                     6880 => "10101101",
                     6881 => "00100101",
                     6882 => "00000111",
                     6883 => "10010101",
                     6884 => "01101110",
                     6885 => "00100000",
                     6886 => "11010101",
                     6887 => "10011011",
                     6888 => "10010101",
                     6889 => "11001111",
                     6890 => "10010101",
                     6891 => "01011000",
                     6892 => "10101001",
                     6893 => "00110010",
                     6894 => "10010101",
                     6895 => "00010110",
                     6896 => "10100000",
                     6897 => "00000001",
                     6898 => "10010100",
                     6899 => "10110110",
                     6900 => "11110110",
                     6901 => "00001111",
                     6902 => "10100110",
                     6903 => "00000111",
                     6904 => "10101001",
                     6905 => "01100111",
                     6906 => "10011101",
                     6907 => "10100001",
                     6908 => "00000110",
                     6909 => "10101001",
                     6910 => "01101000",
                     6911 => "10011101",
                     6912 => "10100010",
                     6913 => "00000110",
                     6914 => "01100000",
                     6915 => "10101101",
                     6916 => "01011101",
                     6917 => "00000111",
                     6918 => "11110000",
                     6919 => "00110110",
                     6920 => "10101001",
                     6921 => "00000000",
                     6922 => "10001101",
                     6923 => "01011101",
                     6924 => "00000111",
                     6925 => "01001100",
                     6926 => "00011011",
                     6927 => "10011011",
                     6928 => "00100000",
                     6929 => "00111000",
                     6930 => "10011011",
                     6931 => "01001100",
                     6932 => "00101110",
                     6933 => "10011011",
                     6934 => "10101001",
                     6935 => "00000000",
                     6936 => "10001101",
                     6937 => "10111100",
                     6938 => "00000110",
                     6939 => "00100000",
                     6940 => "00111000",
                     6941 => "10011011",
                     6942 => "10000100",
                     6943 => "00000111",
                     6944 => "10101001",
                     6945 => "00000000",
                     6946 => "10101100",
                     6947 => "01001110",
                     6948 => "00000111",
                     6949 => "10001000",
                     6950 => "11110000",
                     6951 => "00000010",
                     6952 => "10101001",
                     6953 => "00000101",
                     6954 => "00011000",
                     6955 => "01100101",
                     6956 => "00000111",
                     6957 => "10101000",
                     6958 => "10111001",
                     6959 => "11101101",
                     6960 => "10111101",
                     6961 => "01001000",
                     6962 => "00100000",
                     6963 => "10111101",
                     6964 => "10011011",
                     6965 => "01001100",
                     6966 => "01001000",
                     6967 => "10011010",
                     6968 => "10100101",
                     6969 => "00000000",
                     6970 => "00111000",
                     6971 => "11101001",
                     6972 => "00000000",
                     6973 => "10101000",
                     6974 => "01100000",
                     6975 => "10000111",
                     6976 => "00000000",
                     6977 => "00000000",
                     6978 => "00000000",
                     6979 => "00100000",
                     6980 => "10101110",
                     6981 => "10011011",
                     6982 => "10010000",
                     6983 => "00101101",
                     6984 => "10101101",
                     6985 => "01001110",
                     6986 => "00000111",
                     6987 => "11010000",
                     6988 => "00101000",
                     6989 => "10101110",
                     6990 => "01101010",
                     6991 => "00000100",
                     6992 => "00100000",
                     6993 => "11001101",
                     6994 => "10011011",
                     6995 => "00111000",
                     6996 => "11101001",
                     6997 => "00010000",
                     6998 => "10011101",
                     6999 => "01110001",
                     7000 => "00000100",
                     7001 => "10101101",
                     7002 => "00100101",
                     7003 => "00000111",
                     7004 => "11101001",
                     7005 => "00000000",
                     7006 => "10011101",
                     7007 => "01101011",
                     7008 => "00000100",
                     7009 => "11001000",
                     7010 => "11001000",
                     7011 => "10011000",
                     7012 => "00001010",
                     7013 => "00001010",
                     7014 => "00001010",
                     7015 => "00001010",
                     7016 => "10011101",
                     7017 => "01110111",
                     7018 => "00000100",
                     7019 => "11101000",
                     7020 => "11100000",
                     7021 => "00000101",
                     7022 => "10010000",
                     7023 => "00000010",
                     7024 => "10100010",
                     7025 => "00000000",
                     7026 => "10001110",
                     7027 => "01101010",
                     7028 => "00000100",
                     7029 => "10101110",
                     7030 => "01001110",
                     7031 => "00000111",
                     7032 => "10111101",
                     7033 => "00111111",
                     7034 => "10011011",
                     7035 => "10100010",
                     7036 => "00001000",
                     7037 => "10100000",
                     7038 => "00001111",
                     7039 => "10001100",
                     7040 => "00110101",
                     7041 => "00000111",
                     7042 => "10111100",
                     7043 => "10100001",
                     7044 => "00000110",
                     7045 => "11110000",
                     7046 => "00011000",
                     7047 => "11000000",
                     7048 => "00010111",
                     7049 => "11110000",
                     7050 => "00010111",
                     7051 => "11000000",
                     7052 => "00011010",
                     7053 => "11110000",
                     7054 => "00010011",
                     7055 => "11000000",
                     7056 => "11000000",
                     7057 => "11110000",
                     7058 => "00001100",
                     7059 => "11000000",
                     7060 => "11000000",
                     7061 => "10110000",
                     7062 => "00001011",
                     7063 => "11000000",
                     7064 => "01010100",
                     7065 => "11010000",
                     7066 => "00000100",
                     7067 => "11001001",
                     7068 => "01010000",
                     7069 => "11110000",
                     7070 => "00000011",
                     7071 => "10011101",
                     7072 => "10100001",
                     7073 => "00000110",
                     7074 => "11101000",
                     7075 => "11100000",
                     7076 => "00001101",
                     7077 => "10110000",
                     7078 => "00000110",
                     7079 => "10101100",
                     7080 => "00110101",
                     7081 => "00000111",
                     7082 => "10001000",
                     7083 => "00010000",
                     7084 => "11010010",
                     7085 => "01100000",
                     7086 => "00100000",
                     7087 => "10111101",
                     7088 => "10011011",
                     7089 => "10111101",
                     7090 => "00110000",
                     7091 => "00000111",
                     7092 => "00011000",
                     7093 => "00010000",
                     7094 => "00000101",
                     7095 => "10011000",
                     7096 => "10011101",
                     7097 => "00110000",
                     7098 => "00000111",
                     7099 => "00111000",
                     7100 => "01100000",
                     7101 => "10111100",
                     7102 => "00101101",
                     7103 => "00000111",
                     7104 => "10110001",
                     7105 => "11100111",
                     7106 => "00101001",
                     7107 => "00001111",
                     7108 => "10000101",
                     7109 => "00000111",
                     7110 => "11001000",
                     7111 => "10110001",
                     7112 => "11100111",
                     7113 => "00101001",
                     7114 => "00001111",
                     7115 => "10101000",
                     7116 => "01100000",
                     7117 => "10101101",
                     7118 => "00100110",
                     7119 => "00000111",
                     7120 => "00001010",
                     7121 => "00001010",
                     7122 => "00001010",
                     7123 => "00001010",
                     7124 => "01100000",
                     7125 => "10100101",
                     7126 => "00000111",
                     7127 => "00001010",
                     7128 => "00001010",
                     7129 => "00001010",
                     7130 => "00001010",
                     7131 => "00011000",
                     7132 => "01101001",
                     7133 => "00100000",
                     7134 => "01100000",
                     7135 => "00000000",
                     7136 => "11010000",
                     7137 => "00000101",
                     7138 => "00000101",
                     7139 => "01001000",
                     7140 => "01001010",
                     7141 => "01001010",
                     7142 => "01001010",
                     7143 => "01001010",
                     7144 => "10101000",
                     7145 => "10111001",
                     7146 => "11100001",
                     7147 => "10011011",
                     7148 => "10000101",
                     7149 => "00000111",
                     7150 => "01101000",
                     7151 => "00101001",
                     7152 => "00001111",
                     7153 => "00011000",
                     7154 => "01111001",
                     7155 => "11011111",
                     7156 => "10011011",
                     7157 => "10000101",
                     7158 => "00000110",
                     7159 => "01100000",
                     7160 => "00010010",
                     7161 => "00110110",
                     7162 => "00001110",
                     7163 => "00001110",
                     7164 => "00001110",
                     7165 => "00110010",
                     7166 => "00110010",
                     7167 => "00110010",
                     7168 => "00001010",
                     7169 => "00100110",
                     7170 => "01000000",
                     7171 => "00100000",
                     7172 => "00010011",
                     7173 => "10011100",
                     7174 => "10001101",
                     7175 => "01010000",
                     7176 => "00000111",
                     7177 => "00101001",
                     7178 => "01100000",
                     7179 => "00001010",
                     7180 => "00101010",
                     7181 => "00101010",
                     7182 => "00101010",
                     7183 => "10001101",
                     7184 => "01001110",
                     7185 => "00000111",
                     7186 => "01100000",
                     7187 => "10101100",
                     7188 => "01011111",
                     7189 => "00000111",
                     7190 => "10111001",
                     7191 => "10110100",
                     7192 => "10011100",
                     7193 => "00011000",
                     7194 => "01101101",
                     7195 => "01100000",
                     7196 => "00000111",
                     7197 => "10101000",
                     7198 => "10111001",
                     7199 => "10111100",
                     7200 => "10011100",
                     7201 => "01100000",
                     7202 => "10101101",
                     7203 => "01010000",
                     7204 => "00000111",
                     7205 => "00100000",
                     7206 => "00001001",
                     7207 => "10011100",
                     7208 => "10101000",
                     7209 => "10101101",
                     7210 => "01010000",
                     7211 => "00000111",
                     7212 => "00101001",
                     7213 => "00011111",
                     7214 => "10001101",
                     7215 => "01001111",
                     7216 => "00000111",
                     7217 => "10111001",
                     7218 => "11100000",
                     7219 => "10011100",
                     7220 => "00011000",
                     7221 => "01101101",
                     7222 => "01001111",
                     7223 => "00000111",
                     7224 => "10101000",
                     7225 => "10111001",
                     7226 => "11100100",
                     7227 => "10011100",
                     7228 => "10000101",
                     7229 => "11101001",
                     7230 => "10111001",
                     7231 => "00000110",
                     7232 => "10011101",
                     7233 => "10000101",
                     7234 => "11101010",
                     7235 => "10101100",
                     7236 => "01001110",
                     7237 => "00000111",
                     7238 => "10111001",
                     7239 => "00101000",
                     7240 => "10011101",
                     7241 => "00011000",
                     7242 => "01101101",
                     7243 => "01001111",
                     7244 => "00000111",
                     7245 => "10101000",
                     7246 => "10111001",
                     7247 => "00101100",
                     7248 => "10011101",
                     7249 => "10000101",
                     7250 => "11100111",
                     7251 => "10111001",
                     7252 => "01001110",
                     7253 => "10011101",
                     7254 => "10000101",
                     7255 => "11101000",
                     7256 => "10100000",
                     7257 => "00000000",
                     7258 => "10110001",
                     7259 => "11100111",
                     7260 => "01001000",
                     7261 => "00101001",
                     7262 => "00000111",
                     7263 => "11001001",
                     7264 => "00000100",
                     7265 => "10010000",
                     7266 => "00000101",
                     7267 => "10001101",
                     7268 => "01000100",
                     7269 => "00000111",
                     7270 => "10101001",
                     7271 => "00000000",
                     7272 => "10001101",
                     7273 => "01000001",
                     7274 => "00000111",
                     7275 => "01101000",
                     7276 => "01001000",
                     7277 => "00101001",
                     7278 => "00111000",
                     7279 => "01001010",
                     7280 => "01001010",
                     7281 => "01001010",
                     7282 => "10001101",
                     7283 => "00010000",
                     7284 => "00000111",
                     7285 => "01101000",
                     7286 => "00101001",
                     7287 => "11000000",
                     7288 => "00011000",
                     7289 => "00101010",
                     7290 => "00101010",
                     7291 => "00101010",
                     7292 => "10001101",
                     7293 => "00010101",
                     7294 => "00000111",
                     7295 => "11001000",
                     7296 => "10110001",
                     7297 => "11100111",
                     7298 => "01001000",
                     7299 => "00101001",
                     7300 => "00001111",
                     7301 => "10001101",
                     7302 => "00100111",
                     7303 => "00000111",
                     7304 => "01101000",
                     7305 => "01001000",
                     7306 => "00101001",
                     7307 => "00110000",
                     7308 => "01001010",
                     7309 => "01001010",
                     7310 => "01001010",
                     7311 => "01001010",
                     7312 => "10001101",
                     7313 => "01000010",
                     7314 => "00000111",
                     7315 => "01101000",
                     7316 => "00101001",
                     7317 => "11000000",
                     7318 => "00011000",
                     7319 => "00101010",
                     7320 => "00101010",
                     7321 => "00101010",
                     7322 => "11001001",
                     7323 => "00000011",
                     7324 => "11010000",
                     7325 => "00000101",
                     7326 => "10001101",
                     7327 => "01000011",
                     7328 => "00000111",
                     7329 => "10101001",
                     7330 => "00000000",
                     7331 => "10001101",
                     7332 => "00110011",
                     7333 => "00000111",
                     7334 => "10100101",
                     7335 => "11100111",
                     7336 => "00011000",
                     7337 => "01101001",
                     7338 => "00000010",
                     7339 => "10000101",
                     7340 => "11100111",
                     7341 => "10100101",
                     7342 => "11101000",
                     7343 => "01101001",
                     7344 => "00000000",
                     7345 => "10000101",
                     7346 => "11101000",
                     7347 => "01100000",
                     7348 => "00000000",
                     7349 => "00000101",
                     7350 => "00001010",
                     7351 => "00001110",
                     7352 => "00010011",
                     7353 => "00010111",
                     7354 => "00011011",
                     7355 => "00100000",
                     7356 => "00100101",
                     7357 => "00101001",
                     7358 => "11000000",
                     7359 => "00100110",
                     7360 => "01100000",
                     7361 => "00101000",
                     7362 => "00101001",
                     7363 => "00000001",
                     7364 => "00100111",
                     7365 => "01100010",
                     7366 => "00100100",
                     7367 => "00110101",
                     7368 => "00100000",
                     7369 => "01100011",
                     7370 => "00100010",
                     7371 => "00101001",
                     7372 => "01000001",
                     7373 => "00101100",
                     7374 => "01100001",
                     7375 => "00101010",
                     7376 => "00110001",
                     7377 => "00100110",
                     7378 => "01100010",
                     7379 => "00101110",
                     7380 => "00100011",
                     7381 => "00101101",
                     7382 => "01100000",
                     7383 => "00110011",
                     7384 => "00101001",
                     7385 => "00000001",
                     7386 => "00100111",
                     7387 => "01100100",
                     7388 => "00110000",
                     7389 => "00110010",
                     7390 => "00100001",
                     7391 => "01100101",
                     7392 => "00011111",
                     7393 => "00000110",
                     7394 => "00011100",
                     7395 => "00000000",
                     7396 => "01110000",
                     7397 => "10010111",
                     7398 => "10110000",
                     7399 => "11011111",
                     7400 => "00001010",
                     7401 => "00011111",
                     7402 => "01011001",
                     7403 => "01111110",
                     7404 => "10011011",
                     7405 => "10101001",
                     7406 => "11010000",
                     7407 => "00000001",
                     7408 => "00011111",
                     7409 => "00111100",
                     7410 => "01010001",
                     7411 => "01111011",
                     7412 => "01111100",
                     7413 => "10100000",
                     7414 => "10101001",
                     7415 => "11001110",
                     7416 => "11110001",
                     7417 => "11111010",
                     7418 => "11111011",
                     7419 => "00110101",
                     7420 => "01100000",
                     7421 => "10001110",
                     7422 => "10101010",
                     7423 => "10110011",
                     7424 => "11011000",
                     7425 => "00000101",
                     7426 => "00110011",
                     7427 => "01100000",
                     7428 => "01110001",
                     7429 => "10011011",
                     7430 => "10011101",
                     7431 => "10011101",
                     7432 => "10011101",
                     7433 => "10011101",
                     7434 => "10011110",
                     7435 => "10011110",
                     7436 => "10011110",
                     7437 => "10011110",
                     7438 => "10011110",
                     7439 => "10011110",
                     7440 => "10011110",
                     7441 => "10011111",
                     7442 => "10011111",
                     7443 => "10011111",
                     7444 => "10011111",
                     7445 => "10011111",
                     7446 => "10011111",
                     7447 => "10011111",
                     7448 => "10011111",
                     7449 => "10011111",
                     7450 => "10011111",
                     7451 => "10011111",
                     7452 => "10011111",
                     7453 => "10100000",
                     7454 => "10100000",
                     7455 => "10100000",
                     7456 => "10100000",
                     7457 => "10100000",
                     7458 => "10100000",
                     7459 => "10100001",
                     7460 => "10100001",
                     7461 => "10100001",
                     7462 => "10100001",
                     7463 => "10100001",
                     7464 => "00000000",
                     7465 => "00000011",
                     7466 => "00011001",
                     7467 => "00011100",
                     7468 => "00000110",
                     7469 => "01000101",
                     7470 => "11000000",
                     7471 => "01101011",
                     7472 => "11001110",
                     7473 => "00110111",
                     7474 => "10001010",
                     7475 => "00011001",
                     7476 => "10001110",
                     7477 => "11110011",
                     7478 => "01001000",
                     7479 => "11001101",
                     7480 => "00110010",
                     7481 => "00111011",
                     7482 => "01111010",
                     7483 => "10001111",
                     7484 => "11110110",
                     7485 => "01011011",
                     7486 => "11001110",
                     7487 => "11111111",
                     7488 => "10010010",
                     7489 => "00000101",
                     7490 => "01111110",
                     7491 => "11010111",
                     7492 => "00000010",
                     7493 => "00110101",
                     7494 => "11011000",
                     7495 => "01111001",
                     7496 => "10101111",
                     7497 => "00010000",
                     7498 => "10001111",
                     7499 => "00000010",
                     7500 => "01101111",
                     7501 => "11111010",
                     7502 => "10101110",
                     7503 => "10101110",
                     7504 => "10101110",
                     7505 => "10100100",
                     7506 => "10100100",
                     7507 => "10100101",
                     7508 => "10100101",
                     7509 => "10100110",
                     7510 => "10100110",
                     7511 => "10100110",
                     7512 => "10100111",
                     7513 => "10100111",
                     7514 => "10101000",
                     7515 => "10101000",
                     7516 => "10101000",
                     7517 => "10101000",
                     7518 => "10101000",
                     7519 => "10101001",
                     7520 => "10101001",
                     7521 => "10101001",
                     7522 => "10101010",
                     7523 => "10101011",
                     7524 => "10101011",
                     7525 => "10101011",
                     7526 => "10101100",
                     7527 => "10101100",
                     7528 => "10101100",
                     7529 => "10101101",
                     7530 => "10100001",
                     7531 => "10100010",
                     7532 => "10100010",
                     7533 => "10100011",
                     7534 => "10100011",
                     7535 => "10100011",
                     7536 => "01110110",
                     7537 => "11011101",
                     7538 => "10111011",
                     7539 => "01001100",
                     7540 => "11101010",
                     7541 => "00011101",
                     7542 => "00011011",
                     7543 => "11001100",
                     7544 => "01010110",
                     7545 => "01011101",
                     7546 => "00010110",
                     7547 => "10011101",
                     7548 => "11000110",
                     7549 => "00011101",
                     7550 => "00110110",
                     7551 => "10011101",
                     7552 => "11001001",
                     7553 => "00011101",
                     7554 => "00000100",
                     7555 => "11011011",
                     7556 => "01001001",
                     7557 => "00011101",
                     7558 => "10000100",
                     7559 => "00011011",
                     7560 => "11001001",
                     7561 => "01011101",
                     7562 => "10001000",
                     7563 => "10010101",
                     7564 => "00001111",
                     7565 => "00001000",
                     7566 => "00110000",
                     7567 => "01001100",
                     7568 => "01111000",
                     7569 => "00101101",
                     7570 => "10100110",
                     7571 => "00101000",
                     7572 => "10010000",
                     7573 => "10110101",
                     7574 => "11111111",
                     7575 => "00001111",
                     7576 => "00000011",
                     7577 => "01010110",
                     7578 => "00011011",
                     7579 => "11001001",
                     7580 => "00011011",
                     7581 => "00001111",
                     7582 => "00000111",
                     7583 => "00110110",
                     7584 => "00011011",
                     7585 => "10101010",
                     7586 => "00011011",
                     7587 => "01001000",
                     7588 => "10010101",
                     7589 => "00001111",
                     7590 => "00001010",
                     7591 => "00101010",
                     7592 => "00011011",
                     7593 => "01011011",
                     7594 => "00001100",
                     7595 => "01111000",
                     7596 => "00101101",
                     7597 => "10010000",
                     7598 => "10110101",
                     7599 => "11111111",
                     7600 => "00001011",
                     7601 => "10001100",
                     7602 => "01001011",
                     7603 => "01001100",
                     7604 => "01110111",
                     7605 => "01011111",
                     7606 => "11101011",
                     7607 => "00001100",
                     7608 => "10111101",
                     7609 => "11011011",
                     7610 => "00011001",
                     7611 => "10011101",
                     7612 => "01110101",
                     7613 => "00011101",
                     7614 => "01111101",
                     7615 => "01011011",
                     7616 => "11011001",
                     7617 => "00011101",
                     7618 => "00111101",
                     7619 => "11011101",
                     7620 => "10011001",
                     7621 => "00011101",
                     7622 => "00100110",
                     7623 => "10011101",
                     7624 => "01011010",
                     7625 => "00101011",
                     7626 => "10001010",
                     7627 => "00101100",
                     7628 => "11001010",
                     7629 => "00011011",
                     7630 => "00100000",
                     7631 => "10010101",
                     7632 => "01111011",
                     7633 => "01011100",
                     7634 => "11011011",
                     7635 => "01001100",
                     7636 => "00011011",
                     7637 => "11001100",
                     7638 => "00111011",
                     7639 => "11001100",
                     7640 => "01111000",
                     7641 => "00101101",
                     7642 => "10100110",
                     7643 => "00101000",
                     7644 => "10010000",
                     7645 => "10110101",
                     7646 => "11111111",
                     7647 => "00001011",
                     7648 => "10001100",
                     7649 => "00111011",
                     7650 => "00011101",
                     7651 => "10001011",
                     7652 => "00011101",
                     7653 => "10101011",
                     7654 => "00001100",
                     7655 => "11011011",
                     7656 => "00011101",
                     7657 => "00001111",
                     7658 => "00000011",
                     7659 => "01100101",
                     7660 => "00011101",
                     7661 => "01101011",
                     7662 => "00011011",
                     7663 => "00000101",
                     7664 => "10011101",
                     7665 => "00001011",
                     7666 => "00011011",
                     7667 => "00000101",
                     7668 => "10011011",
                     7669 => "00001011",
                     7670 => "00011101",
                     7671 => "10001011",
                     7672 => "00001100",
                     7673 => "00011011",
                     7674 => "10001100",
                     7675 => "01110000",
                     7676 => "00010101",
                     7677 => "01111011",
                     7678 => "00001100",
                     7679 => "11011011",
                     7680 => "00001100",
                     7681 => "00001111",
                     7682 => "00001000",
                     7683 => "01111000",
                     7684 => "00101101",
                     7685 => "10100110",
                     7686 => "00101000",
                     7687 => "10010000",
                     7688 => "10110101",
                     7689 => "11111111",
                     7690 => "00100111",
                     7691 => "10101001",
                     7692 => "01001011",
                     7693 => "00001100",
                     7694 => "01101000",
                     7695 => "00101001",
                     7696 => "00001111",
                     7697 => "00000110",
                     7698 => "01110111",
                     7699 => "00011011",
                     7700 => "00001111",
                     7701 => "00001011",
                     7702 => "01100000",
                     7703 => "00010101",
                     7704 => "01001011",
                     7705 => "10001100",
                     7706 => "01111000",
                     7707 => "00101101",
                     7708 => "10010000",
                     7709 => "10110101",
                     7710 => "11111111",
                     7711 => "00001111",
                     7712 => "00000011",
                     7713 => "10001110",
                     7714 => "01100101",
                     7715 => "11100001",
                     7716 => "10111011",
                     7717 => "00111000",
                     7718 => "01101101",
                     7719 => "10101000",
                     7720 => "00111110",
                     7721 => "11100101",
                     7722 => "11100111",
                     7723 => "00001111",
                     7724 => "00001000",
                     7725 => "00001011",
                     7726 => "00000010",
                     7727 => "00101011",
                     7728 => "00000010",
                     7729 => "01011110",
                     7730 => "01100101",
                     7731 => "11100001",
                     7732 => "10111011",
                     7733 => "00001110",
                     7734 => "11011011",
                     7735 => "00001110",
                     7736 => "10111011",
                     7737 => "10001110",
                     7738 => "11011011",
                     7739 => "00001110",
                     7740 => "11111110",
                     7741 => "01100101",
                     7742 => "11101100",
                     7743 => "00001111",
                     7744 => "00001101",
                     7745 => "01001110",
                     7746 => "01100101",
                     7747 => "11100001",
                     7748 => "00001111",
                     7749 => "00001110",
                     7750 => "01001110",
                     7751 => "00000010",
                     7752 => "11100000",
                     7753 => "00001111",
                     7754 => "00010000",
                     7755 => "11111110",
                     7756 => "11100101",
                     7757 => "11100001",
                     7758 => "00011011",
                     7759 => "10000101",
                     7760 => "01111011",
                     7761 => "00001100",
                     7762 => "01011011",
                     7763 => "10010101",
                     7764 => "01111000",
                     7765 => "00101101",
                     7766 => "10010000",
                     7767 => "10110101",
                     7768 => "11111111",
                     7769 => "10100101",
                     7770 => "10000110",
                     7771 => "11100100",
                     7772 => "00101000",
                     7773 => "00011000",
                     7774 => "10101000",
                     7775 => "01000101",
                     7776 => "10000011",
                     7777 => "01101001",
                     7778 => "00000011",
                     7779 => "11000110",
                     7780 => "00101001",
                     7781 => "10011011",
                     7782 => "10000011",
                     7783 => "00010110",
                     7784 => "10100100",
                     7785 => "10001000",
                     7786 => "00100100",
                     7787 => "11101001",
                     7788 => "00101000",
                     7789 => "00000101",
                     7790 => "10101000",
                     7791 => "01111011",
                     7792 => "00101000",
                     7793 => "00100100",
                     7794 => "10001111",
                     7795 => "11001000",
                     7796 => "00000011",
                     7797 => "11101000",
                     7798 => "00000011",
                     7799 => "01000110",
                     7800 => "10101000",
                     7801 => "10000101",
                     7802 => "00100100",
                     7803 => "11001000",
                     7804 => "00100100",
                     7805 => "11111111",
                     7806 => "11101011",
                     7807 => "10001110",
                     7808 => "00001111",
                     7809 => "00000011",
                     7810 => "11111011",
                     7811 => "00000101",
                     7812 => "00010111",
                     7813 => "10000101",
                     7814 => "11011011",
                     7815 => "10001110",
                     7816 => "00001111",
                     7817 => "00000111",
                     7818 => "01010111",
                     7819 => "00000101",
                     7820 => "01111011",
                     7821 => "00000101",
                     7822 => "10011011",
                     7823 => "10000000",
                     7824 => "00101011",
                     7825 => "10000101",
                     7826 => "11111011",
                     7827 => "00000101",
                     7828 => "00001111",
                     7829 => "00001011",
                     7830 => "00011011",
                     7831 => "00000101",
                     7832 => "10011011",
                     7833 => "00000101",
                     7834 => "11111111",
                     7835 => "00101110",
                     7836 => "11000010",
                     7837 => "01100110",
                     7838 => "11100010",
                     7839 => "00010001",
                     7840 => "00001111",
                     7841 => "00000111",
                     7842 => "00000010",
                     7843 => "00010001",
                     7844 => "00001111",
                     7845 => "00001100",
                     7846 => "00010010",
                     7847 => "00010001",
                     7848 => "11111111",
                     7849 => "00001110",
                     7850 => "11000010",
                     7851 => "10101000",
                     7852 => "10101011",
                     7853 => "00000000",
                     7854 => "10111011",
                     7855 => "10001110",
                     7856 => "01101011",
                     7857 => "10000010",
                     7858 => "11011110",
                     7859 => "00000000",
                     7860 => "10100000",
                     7861 => "00110011",
                     7862 => "10000110",
                     7863 => "01000011",
                     7864 => "00000110",
                     7865 => "00111110",
                     7866 => "10110100",
                     7867 => "10100000",
                     7868 => "11001011",
                     7869 => "00000010",
                     7870 => "00001111",
                     7871 => "00000111",
                     7872 => "01111110",
                     7873 => "01000010",
                     7874 => "10100110",
                     7875 => "10000011",
                     7876 => "00000010",
                     7877 => "00001111",
                     7878 => "00001010",
                     7879 => "00111011",
                     7880 => "00000010",
                     7881 => "11001011",
                     7882 => "00110111",
                     7883 => "00001111",
                     7884 => "00001100",
                     7885 => "11100011",
                     7886 => "00001110",
                     7887 => "11111111",
                     7888 => "10011011",
                     7889 => "10001110",
                     7890 => "11001010",
                     7891 => "00001110",
                     7892 => "11101110",
                     7893 => "01000010",
                     7894 => "01000100",
                     7895 => "01011011",
                     7896 => "10000110",
                     7897 => "10000000",
                     7898 => "10111000",
                     7899 => "00011011",
                     7900 => "10000000",
                     7901 => "01010000",
                     7902 => "10111010",
                     7903 => "00010000",
                     7904 => "10110111",
                     7905 => "01011011",
                     7906 => "00000000",
                     7907 => "00010111",
                     7908 => "10000101",
                     7909 => "01001011",
                     7910 => "00000101",
                     7911 => "11111110",
                     7912 => "00110100",
                     7913 => "01000000",
                     7914 => "10110111",
                     7915 => "10000110",
                     7916 => "11000110",
                     7917 => "00000110",
                     7918 => "01011011",
                     7919 => "10000000",
                     7920 => "10000011",
                     7921 => "00000000",
                     7922 => "11010000",
                     7923 => "00111000",
                     7924 => "01011011",
                     7925 => "10001110",
                     7926 => "10001010",
                     7927 => "00001110",
                     7928 => "10100110",
                     7929 => "00000000",
                     7930 => "10111011",
                     7931 => "00001110",
                     7932 => "11000101",
                     7933 => "10000000",
                     7934 => "11110011",
                     7935 => "00000000",
                     7936 => "11111111",
                     7937 => "00011110",
                     7938 => "11000010",
                     7939 => "00000000",
                     7940 => "01101011",
                     7941 => "00000110",
                     7942 => "10001011",
                     7943 => "10000110",
                     7944 => "01100011",
                     7945 => "10110111",
                     7946 => "00001111",
                     7947 => "00000101",
                     7948 => "00000011",
                     7949 => "00000110",
                     7950 => "00100011",
                     7951 => "00000110",
                     7952 => "01001011",
                     7953 => "10110111",
                     7954 => "10111011",
                     7955 => "00000000",
                     7956 => "01011011",
                     7957 => "10110111",
                     7958 => "11111011",
                     7959 => "00110111",
                     7960 => "00111011",
                     7961 => "10110111",
                     7962 => "00001111",
                     7963 => "00001011",
                     7964 => "00011011",
                     7965 => "00110111",
                     7966 => "11111111",
                     7967 => "00101011",
                     7968 => "11010111",
                     7969 => "11100011",
                     7970 => "00000011",
                     7971 => "11000010",
                     7972 => "10000110",
                     7973 => "11100010",
                     7974 => "00000110",
                     7975 => "01110110",
                     7976 => "10100101",
                     7977 => "10100011",
                     7978 => "10001111",
                     7979 => "00000011",
                     7980 => "10000110",
                     7981 => "00101011",
                     7982 => "01010111",
                     7983 => "01101000",
                     7984 => "00101000",
                     7985 => "11101001",
                     7986 => "00101000",
                     7987 => "11100101",
                     7988 => "10000011",
                     7989 => "00100100",
                     7990 => "10001111",
                     7991 => "00110110",
                     7992 => "10101000",
                     7993 => "01011011",
                     7994 => "00000011",
                     7995 => "11111111",
                     7996 => "00001111",
                     7997 => "00000010",
                     7998 => "01111000",
                     7999 => "01000000",
                     8000 => "01001000",
                     8001 => "11001110",
                     8002 => "11111000",
                     8003 => "11000011",
                     8004 => "11111000",
                     8005 => "11000011",
                     8006 => "00001111",
                     8007 => "00000111",
                     8008 => "01111011",
                     8009 => "01000011",
                     8010 => "11000110",
                     8011 => "11010000",
                     8012 => "00001111",
                     8013 => "10001010",
                     8014 => "11001000",
                     8015 => "01010000",
                     8016 => "11111111",
                     8017 => "10000101",
                     8018 => "10000110",
                     8019 => "00001011",
                     8020 => "10000000",
                     8021 => "00011011",
                     8022 => "00000000",
                     8023 => "11011011",
                     8024 => "00110111",
                     8025 => "01110111",
                     8026 => "10000000",
                     8027 => "11101011",
                     8028 => "00110111",
                     8029 => "11111110",
                     8030 => "00101011",
                     8031 => "00100000",
                     8032 => "00101011",
                     8033 => "10000000",
                     8034 => "01111011",
                     8035 => "00111000",
                     8036 => "10101011",
                     8037 => "10111000",
                     8038 => "01110111",
                     8039 => "10000110",
                     8040 => "11111110",
                     8041 => "01000010",
                     8042 => "00100000",
                     8043 => "01001001",
                     8044 => "10000110",
                     8045 => "10001011",
                     8046 => "00000110",
                     8047 => "10011011",
                     8048 => "10000000",
                     8049 => "01111011",
                     8050 => "10001110",
                     8051 => "01011011",
                     8052 => "10110111",
                     8053 => "10011011",
                     8054 => "00001110",
                     8055 => "10111011",
                     8056 => "00001110",
                     8057 => "10011011",
                     8058 => "10000000",
                     8059 => "11111111",
                     8060 => "00001011",
                     8061 => "10000000",
                     8062 => "01100000",
                     8063 => "00111000",
                     8064 => "00010000",
                     8065 => "10111000",
                     8066 => "11000000",
                     8067 => "00111011",
                     8068 => "11011011",
                     8069 => "10001110",
                     8070 => "01000000",
                     8071 => "10111000",
                     8072 => "11110000",
                     8073 => "00111000",
                     8074 => "01111011",
                     8075 => "10001110",
                     8076 => "10100000",
                     8077 => "10111000",
                     8078 => "11000000",
                     8079 => "10111000",
                     8080 => "11111011",
                     8081 => "00000000",
                     8082 => "10100000",
                     8083 => "10111000",
                     8084 => "00110000",
                     8085 => "10111011",
                     8086 => "11101110",
                     8087 => "01000010",
                     8088 => "10001000",
                     8089 => "00001111",
                     8090 => "00001011",
                     8091 => "00101011",
                     8092 => "00001110",
                     8093 => "01100111",
                     8094 => "00001110",
                     8095 => "11111111",
                     8096 => "00001010",
                     8097 => "10101010",
                     8098 => "00001110",
                     8099 => "00101000",
                     8100 => "00101010",
                     8101 => "00001110",
                     8102 => "00110001",
                     8103 => "10001000",
                     8104 => "11111111",
                     8105 => "11000111",
                     8106 => "10000011",
                     8107 => "11010111",
                     8108 => "00000011",
                     8109 => "01000010",
                     8110 => "10001111",
                     8111 => "01111010",
                     8112 => "00000011",
                     8113 => "00000101",
                     8114 => "10100100",
                     8115 => "01111000",
                     8116 => "00100100",
                     8117 => "10100110",
                     8118 => "00100101",
                     8119 => "11100100",
                     8120 => "00100101",
                     8121 => "01001011",
                     8122 => "10000011",
                     8123 => "11100011",
                     8124 => "00000011",
                     8125 => "00000101",
                     8126 => "10100100",
                     8127 => "10001001",
                     8128 => "00100100",
                     8129 => "10110101",
                     8130 => "00100100",
                     8131 => "00001001",
                     8132 => "10100100",
                     8133 => "01100101",
                     8134 => "00100100",
                     8135 => "11001001",
                     8136 => "00100100",
                     8137 => "00001111",
                     8138 => "00001000",
                     8139 => "10000101",
                     8140 => "00100101",
                     8141 => "11111111",
                     8142 => "11001101",
                     8143 => "10100101",
                     8144 => "10110101",
                     8145 => "10101000",
                     8146 => "00000111",
                     8147 => "10101000",
                     8148 => "01110110",
                     8149 => "00101000",
                     8150 => "11001100",
                     8151 => "00100101",
                     8152 => "01100101",
                     8153 => "10100100",
                     8154 => "10101001",
                     8155 => "00100100",
                     8156 => "11100101",
                     8157 => "00100100",
                     8158 => "00011001",
                     8159 => "10100100",
                     8160 => "00001111",
                     8161 => "00000111",
                     8162 => "10010101",
                     8163 => "00101000",
                     8164 => "11100110",
                     8165 => "00100100",
                     8166 => "00011001",
                     8167 => "10100100",
                     8168 => "11010111",
                     8169 => "00101001",
                     8170 => "00010110",
                     8171 => "10101001",
                     8172 => "01011000",
                     8173 => "00101001",
                     8174 => "10010111",
                     8175 => "00101001",
                     8176 => "11111111",
                     8177 => "00001111",
                     8178 => "00000010",
                     8179 => "00000010",
                     8180 => "00010001",
                     8181 => "00001111",
                     8182 => "00000111",
                     8183 => "00000010",
                     8184 => "00010001",
                     8185 => "11111111",
                     8186 => "11111111",
                     8187 => "00101011",
                     8188 => "10000010",
                     8189 => "10101011",
                     8190 => "00111000",
                     8191 => "11011110",
                     8192 => "01000010",
                     8193 => "11100010",
                     8194 => "00011011",
                     8195 => "10111000",
                     8196 => "11101011",
                     8197 => "00111011",
                     8198 => "11011011",
                     8199 => "10000000",
                     8200 => "10001011",
                     8201 => "10111000",
                     8202 => "00011011",
                     8203 => "10000010",
                     8204 => "11111011",
                     8205 => "10111000",
                     8206 => "01111011",
                     8207 => "10000000",
                     8208 => "11111011",
                     8209 => "00111100",
                     8210 => "01011011",
                     8211 => "10111100",
                     8212 => "01111011",
                     8213 => "10111000",
                     8214 => "00011011",
                     8215 => "10001110",
                     8216 => "11001011",
                     8217 => "00001110",
                     8218 => "00011011",
                     8219 => "10001110",
                     8220 => "00001111",
                     8221 => "00001101",
                     8222 => "00101011",
                     8223 => "00111011",
                     8224 => "10111011",
                     8225 => "10111000",
                     8226 => "11101011",
                     8227 => "10000010",
                     8228 => "01001011",
                     8229 => "10111000",
                     8230 => "10111011",
                     8231 => "00111000",
                     8232 => "00111011",
                     8233 => "10110111",
                     8234 => "10111011",
                     8235 => "00000010",
                     8236 => "00001111",
                     8237 => "00010011",
                     8238 => "00011011",
                     8239 => "00000000",
                     8240 => "11001011",
                     8241 => "10000000",
                     8242 => "01101011",
                     8243 => "10111100",
                     8244 => "11111111",
                     8245 => "01111011",
                     8246 => "10000000",
                     8247 => "10101110",
                     8248 => "00000000",
                     8249 => "10000000",
                     8250 => "10001011",
                     8251 => "10001110",
                     8252 => "11101000",
                     8253 => "00000101",
                     8254 => "11111001",
                     8255 => "10000110",
                     8256 => "00010111",
                     8257 => "10000110",
                     8258 => "00010110",
                     8259 => "10000101",
                     8260 => "01001110",
                     8261 => "00101011",
                     8262 => "10000000",
                     8263 => "10101011",
                     8264 => "10001110",
                     8265 => "10000111",
                     8266 => "10000101",
                     8267 => "11000011",
                     8268 => "00000101",
                     8269 => "10001011",
                     8270 => "10000010",
                     8271 => "10011011",
                     8272 => "00000010",
                     8273 => "10101011",
                     8274 => "00000010",
                     8275 => "10111011",
                     8276 => "10000110",
                     8277 => "11001011",
                     8278 => "00000110",
                     8279 => "11010011",
                     8280 => "00000011",
                     8281 => "00111011",
                     8282 => "10001110",
                     8283 => "01101011",
                     8284 => "00001110",
                     8285 => "10100111",
                     8286 => "10001110",
                     8287 => "11111111",
                     8288 => "00011001",
                     8289 => "10001110",
                     8290 => "01010010",
                     8291 => "00010001",
                     8292 => "10010011",
                     8293 => "00001110",
                     8294 => "00001111",
                     8295 => "00000011",
                     8296 => "10011011",
                     8297 => "00001110",
                     8298 => "00101011",
                     8299 => "10001110",
                     8300 => "01011011",
                     8301 => "00001110",
                     8302 => "11001011",
                     8303 => "10001110",
                     8304 => "11111011",
                     8305 => "00001110",
                     8306 => "11111011",
                     8307 => "10000010",
                     8308 => "10011011",
                     8309 => "10000010",
                     8310 => "10111011",
                     8311 => "00000010",
                     8312 => "11111110",
                     8313 => "01000010",
                     8314 => "11101000",
                     8315 => "10111011",
                     8316 => "10001110",
                     8317 => "00001111",
                     8318 => "00001010",
                     8319 => "10101011",
                     8320 => "00001110",
                     8321 => "11001011",
                     8322 => "00001110",
                     8323 => "11111001",
                     8324 => "00001110",
                     8325 => "10001000",
                     8326 => "10000110",
                     8327 => "10100110",
                     8328 => "00000110",
                     8329 => "11011011",
                     8330 => "00000010",
                     8331 => "10110110",
                     8332 => "10001110",
                     8333 => "11111111",
                     8334 => "10101011",
                     8335 => "11001110",
                     8336 => "11011110",
                     8337 => "01000010",
                     8338 => "11000000",
                     8339 => "11001011",
                     8340 => "11001110",
                     8341 => "01011011",
                     8342 => "10001110",
                     8343 => "00011011",
                     8344 => "11001110",
                     8345 => "01001011",
                     8346 => "10000101",
                     8347 => "01100111",
                     8348 => "01000101",
                     8349 => "00001111",
                     8350 => "00000111",
                     8351 => "00101011",
                     8352 => "00000000",
                     8353 => "01111011",
                     8354 => "10000101",
                     8355 => "10010111",
                     8356 => "00000101",
                     8357 => "00001111",
                     8358 => "00001010",
                     8359 => "10010010",
                     8360 => "00000010",
                     8361 => "11111111",
                     8362 => "00001010",
                     8363 => "10101010",
                     8364 => "00001110",
                     8365 => "00100100",
                     8366 => "01001010",
                     8367 => "00011110",
                     8368 => "00100011",
                     8369 => "10101010",
                     8370 => "11111111",
                     8371 => "00011011",
                     8372 => "10000000",
                     8373 => "10111011",
                     8374 => "00111000",
                     8375 => "01001011",
                     8376 => "10111100",
                     8377 => "11101011",
                     8378 => "00111011",
                     8379 => "00001111",
                     8380 => "00000100",
                     8381 => "00101011",
                     8382 => "00000000",
                     8383 => "10101011",
                     8384 => "00111000",
                     8385 => "11101011",
                     8386 => "00000000",
                     8387 => "11001011",
                     8388 => "10001110",
                     8389 => "11111011",
                     8390 => "10000000",
                     8391 => "10101011",
                     8392 => "10111000",
                     8393 => "01101011",
                     8394 => "10000000",
                     8395 => "11111011",
                     8396 => "00111100",
                     8397 => "10011011",
                     8398 => "10111011",
                     8399 => "01011011",
                     8400 => "10111100",
                     8401 => "11111011",
                     8402 => "00000000",
                     8403 => "01101011",
                     8404 => "10111000",
                     8405 => "11111011",
                     8406 => "00111000",
                     8407 => "11111111",
                     8408 => "00001011",
                     8409 => "10000110",
                     8410 => "00011010",
                     8411 => "00000110",
                     8412 => "11011011",
                     8413 => "00000110",
                     8414 => "11011110",
                     8415 => "11000010",
                     8416 => "00000010",
                     8417 => "11110000",
                     8418 => "00111011",
                     8419 => "10111011",
                     8420 => "10000000",
                     8421 => "11101011",
                     8422 => "00000110",
                     8423 => "00001011",
                     8424 => "10000110",
                     8425 => "10010011",
                     8426 => "00000110",
                     8427 => "11110000",
                     8428 => "00111001",
                     8429 => "00001111",
                     8430 => "00000110",
                     8431 => "01100000",
                     8432 => "10111000",
                     8433 => "00011011",
                     8434 => "10000110",
                     8435 => "10100000",
                     8436 => "10111001",
                     8437 => "10110111",
                     8438 => "00100111",
                     8439 => "10111101",
                     8440 => "00100111",
                     8441 => "00101011",
                     8442 => "10000011",
                     8443 => "10100001",
                     8444 => "00100110",
                     8445 => "10101001",
                     8446 => "00100110",
                     8447 => "11101110",
                     8448 => "00100101",
                     8449 => "00001011",
                     8450 => "00100111",
                     8451 => "10110100",
                     8452 => "11111111",
                     8453 => "00001111",
                     8454 => "00000010",
                     8455 => "00011110",
                     8456 => "00101111",
                     8457 => "01100000",
                     8458 => "11100000",
                     8459 => "00111010",
                     8460 => "10100101",
                     8461 => "10100111",
                     8462 => "11011011",
                     8463 => "10000000",
                     8464 => "00111011",
                     8465 => "10000010",
                     8466 => "10001011",
                     8467 => "00000010",
                     8468 => "11111110",
                     8469 => "01000010",
                     8470 => "01101000",
                     8471 => "01110000",
                     8472 => "10111011",
                     8473 => "00100101",
                     8474 => "10100111",
                     8475 => "00101100",
                     8476 => "00100111",
                     8477 => "10110010",
                     8478 => "00100110",
                     8479 => "10111001",
                     8480 => "00100110",
                     8481 => "10011011",
                     8482 => "10000000",
                     8483 => "10101000",
                     8484 => "10000010",
                     8485 => "10110101",
                     8486 => "00100111",
                     8487 => "10111100",
                     8488 => "00100111",
                     8489 => "10110000",
                     8490 => "10111011",
                     8491 => "00111011",
                     8492 => "10000010",
                     8493 => "10000111",
                     8494 => "00110100",
                     8495 => "11101110",
                     8496 => "00100101",
                     8497 => "01101011",
                     8498 => "11111111",
                     8499 => "00011110",
                     8500 => "10100101",
                     8501 => "00001010",
                     8502 => "00101110",
                     8503 => "00101000",
                     8504 => "00100111",
                     8505 => "00101110",
                     8506 => "00110011",
                     8507 => "11000111",
                     8508 => "00001111",
                     8509 => "00000011",
                     8510 => "00011110",
                     8511 => "01000000",
                     8512 => "00000111",
                     8513 => "00101110",
                     8514 => "00110000",
                     8515 => "11100111",
                     8516 => "00001111",
                     8517 => "00000101",
                     8518 => "00011110",
                     8519 => "00100100",
                     8520 => "01000100",
                     8521 => "00001111",
                     8522 => "00000111",
                     8523 => "00011110",
                     8524 => "00100010",
                     8525 => "01101010",
                     8526 => "00101110",
                     8527 => "00100011",
                     8528 => "10101011",
                     8529 => "00001111",
                     8530 => "00001001",
                     8531 => "00011110",
                     8532 => "01000001",
                     8533 => "01101000",
                     8534 => "00011110",
                     8535 => "00101010",
                     8536 => "10001010",
                     8537 => "00101110",
                     8538 => "00100011",
                     8539 => "10100010",
                     8540 => "00101110",
                     8541 => "00110010",
                     8542 => "11101010",
                     8543 => "11111111",
                     8544 => "00111011",
                     8545 => "10000111",
                     8546 => "01100110",
                     8547 => "00100111",
                     8548 => "11001100",
                     8549 => "00100111",
                     8550 => "11101110",
                     8551 => "00110001",
                     8552 => "10000111",
                     8553 => "11101110",
                     8554 => "00100011",
                     8555 => "10100111",
                     8556 => "00111011",
                     8557 => "10000111",
                     8558 => "11011011",
                     8559 => "00000111",
                     8560 => "11111111",
                     8561 => "00001111",
                     8562 => "00000001",
                     8563 => "00101110",
                     8564 => "00100101",
                     8565 => "00101011",
                     8566 => "00101110",
                     8567 => "00100101",
                     8568 => "01001011",
                     8569 => "01001110",
                     8570 => "00100101",
                     8571 => "11001011",
                     8572 => "01101011",
                     8573 => "00000111",
                     8574 => "10010111",
                     8575 => "01000111",
                     8576 => "11101001",
                     8577 => "10000111",
                     8578 => "01000111",
                     8579 => "11000111",
                     8580 => "01111010",
                     8581 => "00000111",
                     8582 => "11010110",
                     8583 => "11000111",
                     8584 => "01111000",
                     8585 => "00000111",
                     8586 => "00111000",
                     8587 => "10000111",
                     8588 => "10101011",
                     8589 => "01000111",
                     8590 => "11100011",
                     8591 => "00000111",
                     8592 => "10011011",
                     8593 => "10000111",
                     8594 => "00001111",
                     8595 => "00001001",
                     8596 => "01101000",
                     8597 => "01000111",
                     8598 => "11011011",
                     8599 => "11000111",
                     8600 => "00111011",
                     8601 => "11000111",
                     8602 => "11111111",
                     8603 => "01000111",
                     8604 => "10011011",
                     8605 => "11001011",
                     8606 => "00000111",
                     8607 => "11111010",
                     8608 => "00011101",
                     8609 => "10000110",
                     8610 => "10011011",
                     8611 => "00111010",
                     8612 => "10000111",
                     8613 => "01010110",
                     8614 => "00000111",
                     8615 => "10001000",
                     8616 => "00011011",
                     8617 => "00000111",
                     8618 => "10011101",
                     8619 => "00101110",
                     8620 => "01100101",
                     8621 => "11110000",
                     8622 => "11111111",
                     8623 => "10011011",
                     8624 => "00000111",
                     8625 => "00000101",
                     8626 => "00110010",
                     8627 => "00000110",
                     8628 => "00110011",
                     8629 => "00000111",
                     8630 => "00110100",
                     8631 => "11001110",
                     8632 => "00000011",
                     8633 => "11011100",
                     8634 => "01010001",
                     8635 => "11101110",
                     8636 => "00000111",
                     8637 => "01110011",
                     8638 => "11100000",
                     8639 => "01110100",
                     8640 => "00001010",
                     8641 => "01111110",
                     8642 => "00000110",
                     8643 => "10011110",
                     8644 => "00001010",
                     8645 => "11001110",
                     8646 => "00000110",
                     8647 => "11100100",
                     8648 => "00000000",
                     8649 => "11101000",
                     8650 => "00001010",
                     8651 => "11111110",
                     8652 => "00001010",
                     8653 => "00101110",
                     8654 => "10001001",
                     8655 => "01001110",
                     8656 => "00001011",
                     8657 => "01010100",
                     8658 => "00001010",
                     8659 => "00010100",
                     8660 => "10001010",
                     8661 => "11000100",
                     8662 => "00001010",
                     8663 => "00110100",
                     8664 => "10001010",
                     8665 => "01111110",
                     8666 => "00000110",
                     8667 => "11000111",
                     8668 => "00001010",
                     8669 => "00000001",
                     8670 => "11100000",
                     8671 => "00000010",
                     8672 => "00001010",
                     8673 => "01000111",
                     8674 => "00001010",
                     8675 => "10000001",
                     8676 => "01100000",
                     8677 => "10000010",
                     8678 => "00001010",
                     8679 => "11000111",
                     8680 => "00001010",
                     8681 => "00001110",
                     8682 => "10000111",
                     8683 => "01111110",
                     8684 => "00000010",
                     8685 => "10100111",
                     8686 => "00000010",
                     8687 => "10110011",
                     8688 => "00000010",
                     8689 => "11010111",
                     8690 => "00000010",
                     8691 => "11100011",
                     8692 => "00000010",
                     8693 => "00000111",
                     8694 => "10000010",
                     8695 => "00010011",
                     8696 => "00000010",
                     8697 => "00111110",
                     8698 => "00000110",
                     8699 => "01111110",
                     8700 => "00000010",
                     8701 => "10101110",
                     8702 => "00000111",
                     8703 => "11111110",
                     8704 => "00001010",
                     8705 => "00001101",
                     8706 => "11000100",
                     8707 => "11001101",
                     8708 => "01000011",
                     8709 => "11001110",
                     8710 => "00001001",
                     8711 => "11011110",
                     8712 => "00001011",
                     8713 => "11011101",
                     8714 => "01000010",
                     8715 => "11111110",
                     8716 => "00000010",
                     8717 => "01011101",
                     8718 => "11000111",
                     8719 => "11111101",
                     8720 => "01011011",
                     8721 => "00000111",
                     8722 => "00000101",
                     8723 => "00110010",
                     8724 => "00000110",
                     8725 => "00110011",
                     8726 => "00000111",
                     8727 => "00110100",
                     8728 => "01011110",
                     8729 => "00001010",
                     8730 => "01101000",
                     8731 => "01100100",
                     8732 => "10011000",
                     8733 => "01100100",
                     8734 => "10101000",
                     8735 => "01100100",
                     8736 => "11001110",
                     8737 => "00000110",
                     8738 => "11111110",
                     8739 => "00000010",
                     8740 => "00001101",
                     8741 => "00000001",
                     8742 => "00011110",
                     8743 => "00001110",
                     8744 => "01111110",
                     8745 => "00000010",
                     8746 => "10010100",
                     8747 => "01100011",
                     8748 => "10110100",
                     8749 => "01100011",
                     8750 => "11010100",
                     8751 => "01100011",
                     8752 => "11110100",
                     8753 => "01100011",
                     8754 => "00010100",
                     8755 => "11100011",
                     8756 => "00101110",
                     8757 => "00001110",
                     8758 => "01011110",
                     8759 => "00000010",
                     8760 => "01100100",
                     8761 => "00110101",
                     8762 => "10001000",
                     8763 => "01110010",
                     8764 => "10111110",
                     8765 => "00001110",
                     8766 => "00001101",
                     8767 => "00000100",
                     8768 => "10101110",
                     8769 => "00000010",
                     8770 => "11001110",
                     8771 => "00001000",
                     8772 => "11001101",
                     8773 => "01001011",
                     8774 => "11111110",
                     8775 => "00000010",
                     8776 => "00001101",
                     8777 => "00000101",
                     8778 => "01101000",
                     8779 => "00110001",
                     8780 => "01111110",
                     8781 => "00001010",
                     8782 => "10010110",
                     8783 => "00110001",
                     8784 => "10101001",
                     8785 => "01100011",
                     8786 => "10101000",
                     8787 => "00110011",
                     8788 => "11010101",
                     8789 => "00110000",
                     8790 => "11101110",
                     8791 => "00000010",
                     8792 => "11100110",
                     8793 => "01100010",
                     8794 => "11110100",
                     8795 => "01100001",
                     8796 => "00000100",
                     8797 => "10110001",
                     8798 => "00001000",
                     8799 => "00111111",
                     8800 => "01000100",
                     8801 => "00110011",
                     8802 => "10010100",
                     8803 => "01100011",
                     8804 => "10100100",
                     8805 => "00110001",
                     8806 => "11100100",
                     8807 => "00110001",
                     8808 => "00000100",
                     8809 => "10111111",
                     8810 => "00001000",
                     8811 => "00111111",
                     8812 => "00000100",
                     8813 => "10111111",
                     8814 => "00001000",
                     8815 => "00111111",
                     8816 => "11001101",
                     8817 => "01001011",
                     8818 => "00000011",
                     8819 => "11100100",
                     8820 => "00001110",
                     8821 => "00000011",
                     8822 => "00101110",
                     8823 => "00000001",
                     8824 => "01111110",
                     8825 => "00000110",
                     8826 => "10111110",
                     8827 => "00000010",
                     8828 => "11011110",
                     8829 => "00000110",
                     8830 => "11111110",
                     8831 => "00001010",
                     8832 => "00001101",
                     8833 => "11000100",
                     8834 => "11001101",
                     8835 => "01000011",
                     8836 => "11001110",
                     8837 => "00001001",
                     8838 => "11011110",
                     8839 => "00001011",
                     8840 => "11011101",
                     8841 => "01000010",
                     8842 => "11111110",
                     8843 => "00000010",
                     8844 => "01011101",
                     8845 => "11000111",
                     8846 => "11111101",
                     8847 => "10011011",
                     8848 => "00000111",
                     8849 => "00000101",
                     8850 => "00110010",
                     8851 => "00000110",
                     8852 => "00110011",
                     8853 => "00000111",
                     8854 => "00110100",
                     8855 => "11111110",
                     8856 => "00000000",
                     8857 => "00100111",
                     8858 => "10110001",
                     8859 => "01100101",
                     8860 => "00110010",
                     8861 => "01110101",
                     8862 => "00001010",
                     8863 => "01110001",
                     8864 => "00000000",
                     8865 => "10110111",
                     8866 => "00110001",
                     8867 => "00001000",
                     8868 => "11100100",
                     8869 => "00011000",
                     8870 => "01100100",
                     8871 => "00011110",
                     8872 => "00000100",
                     8873 => "01010111",
                     8874 => "00111011",
                     8875 => "10111011",
                     8876 => "00001010",
                     8877 => "00010111",
                     8878 => "10001010",
                     8879 => "00100111",
                     8880 => "00111010",
                     8881 => "01110011",
                     8882 => "00001010",
                     8883 => "01111011",
                     8884 => "00001010",
                     8885 => "11010111",
                     8886 => "00001010",
                     8887 => "11100111",
                     8888 => "00111010",
                     8889 => "00111011",
                     8890 => "10001010",
                     8891 => "10010111",
                     8892 => "00001010",
                     8893 => "11111110",
                     8894 => "00001000",
                     8895 => "00100100",
                     8896 => "10001010",
                     8897 => "00101110",
                     8898 => "00000000",
                     8899 => "00111110",
                     8900 => "01000000",
                     8901 => "00111000",
                     8902 => "01100100",
                     8903 => "01101111",
                     8904 => "00000000",
                     8905 => "10011111",
                     8906 => "00000000",
                     8907 => "10111110",
                     8908 => "01000011",
                     8909 => "11001000",
                     8910 => "00001010",
                     8911 => "11001001",
                     8912 => "01100011",
                     8913 => "11001110",
                     8914 => "00000111",
                     8915 => "11111110",
                     8916 => "00000111",
                     8917 => "00101110",
                     8918 => "10000001",
                     8919 => "01100110",
                     8920 => "01000010",
                     8921 => "01101010",
                     8922 => "01000010",
                     8923 => "01111001",
                     8924 => "00001010",
                     8925 => "10111110",
                     8926 => "00000000",
                     8927 => "11001000",
                     8928 => "01100100",
                     8929 => "11111000",
                     8930 => "01100100",
                     8931 => "00001000",
                     8932 => "11100100",
                     8933 => "00101110",
                     8934 => "00000111",
                     8935 => "01111110",
                     8936 => "00000011",
                     8937 => "10011110",
                     8938 => "00000111",
                     8939 => "10111110",
                     8940 => "00000011",
                     8941 => "11011110",
                     8942 => "00000111",
                     8943 => "11111110",
                     8944 => "00001010",
                     8945 => "00000011",
                     8946 => "10100101",
                     8947 => "00001101",
                     8948 => "01000100",
                     8949 => "11001101",
                     8950 => "01000011",
                     8951 => "11001110",
                     8952 => "00001001",
                     8953 => "11011101",
                     8954 => "01000010",
                     8955 => "11011110",
                     8956 => "00001011",
                     8957 => "11111110",
                     8958 => "00000010",
                     8959 => "01011101",
                     8960 => "11000111",
                     8961 => "11111101",
                     8962 => "10011011",
                     8963 => "00000111",
                     8964 => "00000101",
                     8965 => "00110010",
                     8966 => "00000110",
                     8967 => "00110011",
                     8968 => "00000111",
                     8969 => "00110100",
                     8970 => "11111110",
                     8971 => "00000110",
                     8972 => "00001100",
                     8973 => "10000001",
                     8974 => "00111001",
                     8975 => "00001010",
                     8976 => "01011100",
                     8977 => "00000001",
                     8978 => "10001001",
                     8979 => "00001010",
                     8980 => "10101100",
                     8981 => "00000001",
                     8982 => "11011001",
                     8983 => "00001010",
                     8984 => "11111100",
                     8985 => "00000001",
                     8986 => "00101110",
                     8987 => "10000011",
                     8988 => "10100111",
                     8989 => "00000001",
                     8990 => "10110111",
                     8991 => "00000000",
                     8992 => "11000111",
                     8993 => "00000001",
                     8994 => "11011110",
                     8995 => "00001010",
                     8996 => "11111110",
                     8997 => "00000010",
                     8998 => "01001110",
                     8999 => "10000011",
                     9000 => "01011010",
                     9001 => "00110010",
                     9002 => "01100011",
                     9003 => "00001010",
                     9004 => "01101001",
                     9005 => "00001010",
                     9006 => "01111110",
                     9007 => "00000010",
                     9008 => "11101110",
                     9009 => "00000011",
                     9010 => "11111010",
                     9011 => "00110010",
                     9012 => "00000011",
                     9013 => "10001010",
                     9014 => "00001001",
                     9015 => "00001010",
                     9016 => "00011110",
                     9017 => "00000010",
                     9018 => "11101110",
                     9019 => "00000011",
                     9020 => "11111010",
                     9021 => "00110010",
                     9022 => "00000011",
                     9023 => "10001010",
                     9024 => "00001001",
                     9025 => "00001010",
                     9026 => "00010100",
                     9027 => "01000010",
                     9028 => "00011110",
                     9029 => "00000010",
                     9030 => "01111110",
                     9031 => "00001010",
                     9032 => "10011110",
                     9033 => "00000111",
                     9034 => "11111110",
                     9035 => "00001010",
                     9036 => "00101110",
                     9037 => "10000110",
                     9038 => "01011110",
                     9039 => "00001010",
                     9040 => "10001110",
                     9041 => "00000110",
                     9042 => "10111110",
                     9043 => "00001010",
                     9044 => "11101110",
                     9045 => "00000111",
                     9046 => "00111110",
                     9047 => "10000011",
                     9048 => "01011110",
                     9049 => "00000111",
                     9050 => "11111110",
                     9051 => "00001010",
                     9052 => "00001101",
                     9053 => "11000100",
                     9054 => "01000001",
                     9055 => "01010010",
                     9056 => "01010001",
                     9057 => "01010010",
                     9058 => "11001101",
                     9059 => "01000011",
                     9060 => "11001110",
                     9061 => "00001001",
                     9062 => "11011110",
                     9063 => "00001011",
                     9064 => "11011101",
                     9065 => "01000010",
                     9066 => "11111110",
                     9067 => "00000010",
                     9068 => "01011101",
                     9069 => "11000111",
                     9070 => "11111101",
                     9071 => "01011011",
                     9072 => "00000111",
                     9073 => "00000101",
                     9074 => "00110010",
                     9075 => "00000110",
                     9076 => "00110011",
                     9077 => "00000111",
                     9078 => "00110100",
                     9079 => "11111110",
                     9080 => "00001010",
                     9081 => "10101110",
                     9082 => "10000110",
                     9083 => "10111110",
                     9084 => "00000111",
                     9085 => "11111110",
                     9086 => "00000010",
                     9087 => "00001101",
                     9088 => "00000010",
                     9089 => "00100111",
                     9090 => "00110010",
                     9091 => "01000110",
                     9092 => "01100001",
                     9093 => "01010101",
                     9094 => "01100010",
                     9095 => "01011110",
                     9096 => "00001110",
                     9097 => "00011110",
                     9098 => "10000010",
                     9099 => "01101000",
                     9100 => "00111100",
                     9101 => "01110100",
                     9102 => "00111010",
                     9103 => "01111101",
                     9104 => "01001011",
                     9105 => "01011110",
                     9106 => "10001110",
                     9107 => "01111101",
                     9108 => "01001011",
                     9109 => "01111110",
                     9110 => "10000010",
                     9111 => "10000100",
                     9112 => "01100010",
                     9113 => "10010100",
                     9114 => "01100001",
                     9115 => "10100100",
                     9116 => "00110001",
                     9117 => "10111101",
                     9118 => "01001011",
                     9119 => "11001110",
                     9120 => "00000110",
                     9121 => "11111110",
                     9122 => "00000010",
                     9123 => "00001101",
                     9124 => "00000110",
                     9125 => "00110100",
                     9126 => "00110001",
                     9127 => "00111110",
                     9128 => "00001010",
                     9129 => "01100100",
                     9130 => "00110010",
                     9131 => "01110101",
                     9132 => "00001010",
                     9133 => "01111011",
                     9134 => "01100001",
                     9135 => "10100100",
                     9136 => "00110011",
                     9137 => "10101110",
                     9138 => "00000010",
                     9139 => "11011110",
                     9140 => "00001110",
                     9141 => "00111110",
                     9142 => "10000010",
                     9143 => "01100100",
                     9144 => "00110010",
                     9145 => "01111000",
                     9146 => "00110010",
                     9147 => "10110100",
                     9148 => "00110110",
                     9149 => "11001000",
                     9150 => "00110110",
                     9151 => "11011101",
                     9152 => "01001011",
                     9153 => "01000100",
                     9154 => "10110010",
                     9155 => "01011000",
                     9156 => "00110010",
                     9157 => "10010100",
                     9158 => "01100011",
                     9159 => "10100100",
                     9160 => "00111110",
                     9161 => "10111010",
                     9162 => "00110000",
                     9163 => "11001001",
                     9164 => "01100001",
                     9165 => "11001110",
                     9166 => "00000110",
                     9167 => "11011101",
                     9168 => "01001011",
                     9169 => "11001110",
                     9170 => "10000110",
                     9171 => "11011101",
                     9172 => "01001011",
                     9173 => "11111110",
                     9174 => "00000010",
                     9175 => "00101110",
                     9176 => "10000110",
                     9177 => "01011110",
                     9178 => "00000010",
                     9179 => "01111110",
                     9180 => "00000110",
                     9181 => "11111110",
                     9182 => "00000010",
                     9183 => "00011110",
                     9184 => "10000110",
                     9185 => "00111110",
                     9186 => "00000010",
                     9187 => "01011110",
                     9188 => "00000110",
                     9189 => "01111110",
                     9190 => "00000010",
                     9191 => "10011110",
                     9192 => "00000110",
                     9193 => "11111110",
                     9194 => "00001010",
                     9195 => "00001101",
                     9196 => "11000100",
                     9197 => "11001101",
                     9198 => "01000011",
                     9199 => "11001110",
                     9200 => "00001001",
                     9201 => "11011110",
                     9202 => "00001011",
                     9203 => "11011101",
                     9204 => "01000010",
                     9205 => "11111110",
                     9206 => "00000010",
                     9207 => "01011101",
                     9208 => "11000111",
                     9209 => "11111101",
                     9210 => "01011011",
                     9211 => "00000110",
                     9212 => "00000101",
                     9213 => "00110010",
                     9214 => "00000110",
                     9215 => "00110011",
                     9216 => "00000111",
                     9217 => "00110100",
                     9218 => "01011110",
                     9219 => "00001010",
                     9220 => "10101110",
                     9221 => "00000010",
                     9222 => "00001101",
                     9223 => "00000001",
                     9224 => "00111001",
                     9225 => "01110011",
                     9226 => "00001101",
                     9227 => "00000011",
                     9228 => "00111001",
                     9229 => "01111011",
                     9230 => "01001101",
                     9231 => "01001011",
                     9232 => "11011110",
                     9233 => "00000110",
                     9234 => "00011110",
                     9235 => "10001010",
                     9236 => "10101110",
                     9237 => "00000110",
                     9238 => "11000100",
                     9239 => "00110011",
                     9240 => "00010110",
                     9241 => "11111110",
                     9242 => "10100101",
                     9243 => "01110111",
                     9244 => "11111110",
                     9245 => "00000010",
                     9246 => "11111110",
                     9247 => "10000010",
                     9248 => "00001101",
                     9249 => "00000111",
                     9250 => "00111001",
                     9251 => "01110011",
                     9252 => "10101000",
                     9253 => "01110100",
                     9254 => "11101101",
                     9255 => "01001011",
                     9256 => "01001001",
                     9257 => "11111011",
                     9258 => "11101000",
                     9259 => "01110100",
                     9260 => "11111110",
                     9261 => "00001010",
                     9262 => "00101110",
                     9263 => "10000010",
                     9264 => "01100111",
                     9265 => "00000010",
                     9266 => "10000100",
                     9267 => "01111010",
                     9268 => "10000111",
                     9269 => "00110001",
                     9270 => "00001101",
                     9271 => "00001011",
                     9272 => "11111110",
                     9273 => "00000010",
                     9274 => "00001101",
                     9275 => "00001100",
                     9276 => "00111001",
                     9277 => "01110011",
                     9278 => "01011110",
                     9279 => "00000110",
                     9280 => "11000110",
                     9281 => "01110110",
                     9282 => "01000101",
                     9283 => "11111111",
                     9284 => "10111110",
                     9285 => "00001010",
                     9286 => "11011101",
                     9287 => "01001000",
                     9288 => "11111110",
                     9289 => "00000110",
                     9290 => "00111101",
                     9291 => "11001011",
                     9292 => "01000110",
                     9293 => "01111110",
                     9294 => "10101101",
                     9295 => "01001010",
                     9296 => "11111110",
                     9297 => "10000010",
                     9298 => "00111001",
                     9299 => "11110011",
                     9300 => "10101001",
                     9301 => "01111011",
                     9302 => "01001110",
                     9303 => "10001010",
                     9304 => "10011110",
                     9305 => "00000111",
                     9306 => "11111110",
                     9307 => "00001010",
                     9308 => "00001101",
                     9309 => "11000100",
                     9310 => "11001101",
                     9311 => "01000011",
                     9312 => "11001110",
                     9313 => "00001001",
                     9314 => "11011110",
                     9315 => "00001011",
                     9316 => "11011101",
                     9317 => "01000010",
                     9318 => "11111110",
                     9319 => "00000010",
                     9320 => "01011101",
                     9321 => "11000111",
                     9322 => "11111101",
                     9323 => "10010100",
                     9324 => "00010001",
                     9325 => "00001111",
                     9326 => "00100110",
                     9327 => "11111110",
                     9328 => "00010000",
                     9329 => "00101000",
                     9330 => "10010100",
                     9331 => "01100101",
                     9332 => "00010101",
                     9333 => "11101011",
                     9334 => "00010010",
                     9335 => "11111010",
                     9336 => "01000001",
                     9337 => "01001010",
                     9338 => "10010110",
                     9339 => "01010100",
                     9340 => "01000000",
                     9341 => "10100100",
                     9342 => "01000010",
                     9343 => "10110111",
                     9344 => "00010011",
                     9345 => "11101001",
                     9346 => "00011001",
                     9347 => "11110101",
                     9348 => "00010101",
                     9349 => "00010001",
                     9350 => "10000000",
                     9351 => "01000111",
                     9352 => "01000010",
                     9353 => "01110001",
                     9354 => "00010011",
                     9355 => "10000000",
                     9356 => "01000001",
                     9357 => "00010101",
                     9358 => "10010010",
                     9359 => "00011011",
                     9360 => "00011111",
                     9361 => "00100100",
                     9362 => "01000000",
                     9363 => "01010101",
                     9364 => "00010010",
                     9365 => "01100100",
                     9366 => "01000000",
                     9367 => "10010101",
                     9368 => "00010010",
                     9369 => "10100100",
                     9370 => "01000000",
                     9371 => "11010010",
                     9372 => "00010010",
                     9373 => "11100001",
                     9374 => "01000000",
                     9375 => "00010011",
                     9376 => "11000000",
                     9377 => "00101100",
                     9378 => "00010111",
                     9379 => "00101111",
                     9380 => "00010010",
                     9381 => "01001001",
                     9382 => "00010011",
                     9383 => "10000011",
                     9384 => "01000000",
                     9385 => "10011111",
                     9386 => "00010100",
                     9387 => "10100011",
                     9388 => "01000000",
                     9389 => "00010111",
                     9390 => "10010010",
                     9391 => "10000011",
                     9392 => "00010011",
                     9393 => "10010010",
                     9394 => "01000001",
                     9395 => "10111001",
                     9396 => "00010100",
                     9397 => "11000101",
                     9398 => "00010010",
                     9399 => "11001000",
                     9400 => "01000000",
                     9401 => "11010100",
                     9402 => "01000000",
                     9403 => "01001011",
                     9404 => "10010010",
                     9405 => "01111000",
                     9406 => "00011011",
                     9407 => "10011100",
                     9408 => "10010100",
                     9409 => "10011111",
                     9410 => "00010001",
                     9411 => "11011111",
                     9412 => "00010100",
                     9413 => "11111110",
                     9414 => "00010001",
                     9415 => "01111101",
                     9416 => "11000001",
                     9417 => "10011110",
                     9418 => "01000010",
                     9419 => "11001111",
                     9420 => "00100000",
                     9421 => "11111101",
                     9422 => "10010000",
                     9423 => "10110001",
                     9424 => "00001111",
                     9425 => "00100110",
                     9426 => "00101001",
                     9427 => "10010001",
                     9428 => "01111110",
                     9429 => "01000010",
                     9430 => "11111110",
                     9431 => "01000000",
                     9432 => "00101000",
                     9433 => "10010010",
                     9434 => "01001110",
                     9435 => "01000010",
                     9436 => "00101110",
                     9437 => "11000000",
                     9438 => "01010111",
                     9439 => "01110011",
                     9440 => "11000011",
                     9441 => "00100101",
                     9442 => "11000111",
                     9443 => "00100111",
                     9444 => "00100011",
                     9445 => "10000100",
                     9446 => "00110011",
                     9447 => "00100000",
                     9448 => "01011100",
                     9449 => "00000001",
                     9450 => "01110111",
                     9451 => "01100011",
                     9452 => "10001000",
                     9453 => "01100010",
                     9454 => "10011001",
                     9455 => "01100001",
                     9456 => "10101010",
                     9457 => "01100000",
                     9458 => "10111100",
                     9459 => "00000001",
                     9460 => "11101110",
                     9461 => "01000010",
                     9462 => "01001110",
                     9463 => "11000000",
                     9464 => "01101001",
                     9465 => "00010001",
                     9466 => "01111110",
                     9467 => "01000010",
                     9468 => "11011110",
                     9469 => "01000000",
                     9470 => "11111000",
                     9471 => "01100010",
                     9472 => "00001110",
                     9473 => "11000010",
                     9474 => "10101110",
                     9475 => "01000000",
                     9476 => "11010111",
                     9477 => "01100011",
                     9478 => "11100111",
                     9479 => "01100011",
                     9480 => "00110011",
                     9481 => "10100111",
                     9482 => "00110111",
                     9483 => "00100111",
                     9484 => "01000011",
                     9485 => "00000100",
                     9486 => "11001100",
                     9487 => "00000001",
                     9488 => "11100111",
                     9489 => "01110011",
                     9490 => "00001100",
                     9491 => "10000001",
                     9492 => "00111110",
                     9493 => "01000010",
                     9494 => "00001101",
                     9495 => "00001010",
                     9496 => "01011110",
                     9497 => "01000000",
                     9498 => "10001000",
                     9499 => "01110010",
                     9500 => "10111110",
                     9501 => "01000010",
                     9502 => "11100111",
                     9503 => "10000111",
                     9504 => "11111110",
                     9505 => "01000000",
                     9506 => "00111001",
                     9507 => "11100001",
                     9508 => "01001110",
                     9509 => "00000000",
                     9510 => "01101001",
                     9511 => "01100000",
                     9512 => "10000111",
                     9513 => "01100000",
                     9514 => "10100101",
                     9515 => "01100000",
                     9516 => "11000011",
                     9517 => "00110001",
                     9518 => "11111110",
                     9519 => "00110001",
                     9520 => "01101101",
                     9521 => "11000001",
                     9522 => "10111110",
                     9523 => "01000010",
                     9524 => "11101111",
                     9525 => "00100000",
                     9526 => "11111101",
                     9527 => "01010010",
                     9528 => "00100001",
                     9529 => "00001111",
                     9530 => "00100000",
                     9531 => "01101110",
                     9532 => "01000000",
                     9533 => "01011000",
                     9534 => "11110010",
                     9535 => "10010011",
                     9536 => "00000001",
                     9537 => "10010111",
                     9538 => "00000000",
                     9539 => "00001100",
                     9540 => "10000001",
                     9541 => "10010111",
                     9542 => "01000000",
                     9543 => "10100110",
                     9544 => "01000001",
                     9545 => "11000111",
                     9546 => "01000000",
                     9547 => "00001101",
                     9548 => "00000100",
                     9549 => "00000011",
                     9550 => "00000001",
                     9551 => "00000111",
                     9552 => "00000001",
                     9553 => "00100011",
                     9554 => "00000001",
                     9555 => "00100111",
                     9556 => "00000001",
                     9557 => "11101100",
                     9558 => "00000011",
                     9559 => "10101100",
                     9560 => "11110011",
                     9561 => "11000011",
                     9562 => "00000011",
                     9563 => "01111000",
                     9564 => "11100010",
                     9565 => "10010100",
                     9566 => "01000011",
                     9567 => "01000111",
                     9568 => "11110011",
                     9569 => "01110100",
                     9570 => "01000011",
                     9571 => "01000111",
                     9572 => "11111011",
                     9573 => "01110100",
                     9574 => "01000011",
                     9575 => "00101100",
                     9576 => "11110001",
                     9577 => "01001100",
                     9578 => "01100011",
                     9579 => "01000111",
                     9580 => "00000000",
                     9581 => "01010111",
                     9582 => "00100001",
                     9583 => "01011100",
                     9584 => "00000001",
                     9585 => "01111100",
                     9586 => "01110010",
                     9587 => "00111001",
                     9588 => "11110001",
                     9589 => "11101100",
                     9590 => "00000010",
                     9591 => "01001100",
                     9592 => "10000001",
                     9593 => "11011000",
                     9594 => "01100010",
                     9595 => "11101100",
                     9596 => "00000001",
                     9597 => "00001101",
                     9598 => "00001101",
                     9599 => "00001111",
                     9600 => "00111000",
                     9601 => "11000111",
                     9602 => "00000111",
                     9603 => "11101101",
                     9604 => "01001010",
                     9605 => "00011101",
                     9606 => "11000001",
                     9607 => "01011111",
                     9608 => "00100110",
                     9609 => "11111101",
                     9610 => "01010100",
                     9611 => "00100001",
                     9612 => "00001111",
                     9613 => "00100110",
                     9614 => "10100111",
                     9615 => "00100010",
                     9616 => "00110111",
                     9617 => "11111011",
                     9618 => "01110011",
                     9619 => "00100000",
                     9620 => "10000011",
                     9621 => "00000111",
                     9622 => "10000111",
                     9623 => "00000010",
                     9624 => "10010011",
                     9625 => "00100000",
                     9626 => "11000111",
                     9627 => "01110011",
                     9628 => "00000100",
                     9629 => "11110001",
                     9630 => "00000110",
                     9631 => "00110001",
                     9632 => "00111001",
                     9633 => "01110001",
                     9634 => "01011001",
                     9635 => "01110001",
                     9636 => "11100111",
                     9637 => "01110011",
                     9638 => "00110111",
                     9639 => "10100000",
                     9640 => "01000111",
                     9641 => "00000100",
                     9642 => "10000110",
                     9643 => "01111100",
                     9644 => "11100101",
                     9645 => "01110001",
                     9646 => "11100111",
                     9647 => "00110001",
                     9648 => "00110011",
                     9649 => "10100100",
                     9650 => "00111001",
                     9651 => "01110001",
                     9652 => "10101001",
                     9653 => "01110001",
                     9654 => "11010011",
                     9655 => "00100011",
                     9656 => "00001000",
                     9657 => "11110010",
                     9658 => "00010011",
                     9659 => "00000101",
                     9660 => "00100111",
                     9661 => "00000010",
                     9662 => "01001001",
                     9663 => "01110001",
                     9664 => "01110101",
                     9665 => "01110101",
                     9666 => "11101000",
                     9667 => "01110010",
                     9668 => "01100111",
                     9669 => "11110011",
                     9670 => "10011001",
                     9671 => "01110001",
                     9672 => "11100111",
                     9673 => "00100000",
                     9674 => "11110100",
                     9675 => "01110010",
                     9676 => "11110111",
                     9677 => "00110001",
                     9678 => "00010111",
                     9679 => "10100000",
                     9680 => "00110011",
                     9681 => "00100000",
                     9682 => "00111001",
                     9683 => "01110001",
                     9684 => "01110011",
                     9685 => "00101000",
                     9686 => "10111100",
                     9687 => "00000101",
                     9688 => "00111001",
                     9689 => "11110001",
                     9690 => "01111001",
                     9691 => "01110001",
                     9692 => "10100110",
                     9693 => "00100001",
                     9694 => "11000011",
                     9695 => "00000110",
                     9696 => "11010011",
                     9697 => "00100000",
                     9698 => "11011100",
                     9699 => "00000000",
                     9700 => "11111100",
                     9701 => "00000000",
                     9702 => "00000111",
                     9703 => "10100010",
                     9704 => "00010011",
                     9705 => "00100001",
                     9706 => "01011111",
                     9707 => "00110010",
                     9708 => "10001100",
                     9709 => "00000000",
                     9710 => "10011000",
                     9711 => "01111010",
                     9712 => "11000111",
                     9713 => "01100011",
                     9714 => "11011001",
                     9715 => "01100001",
                     9716 => "00000011",
                     9717 => "10100010",
                     9718 => "00000111",
                     9719 => "00100010",
                     9720 => "01110100",
                     9721 => "01110010",
                     9722 => "01110111",
                     9723 => "00110001",
                     9724 => "11100111",
                     9725 => "01110011",
                     9726 => "00111001",
                     9727 => "11110001",
                     9728 => "01011000",
                     9729 => "01110010",
                     9730 => "01110111",
                     9731 => "01110011",
                     9732 => "11011000",
                     9733 => "01110010",
                     9734 => "01111111",
                     9735 => "10110001",
                     9736 => "10010111",
                     9737 => "01110011",
                     9738 => "10110110",
                     9739 => "01100100",
                     9740 => "11000101",
                     9741 => "01100101",
                     9742 => "11010100",
                     9743 => "01100110",
                     9744 => "11100011",
                     9745 => "01100111",
                     9746 => "11110011",
                     9747 => "01100111",
                     9748 => "10001101",
                     9749 => "11000001",
                     9750 => "11001111",
                     9751 => "00100110",
                     9752 => "11111101",
                     9753 => "01010010",
                     9754 => "00110001",
                     9755 => "00001111",
                     9756 => "00100000",
                     9757 => "01101110",
                     9758 => "01100110",
                     9759 => "00000111",
                     9760 => "10000001",
                     9761 => "00110110",
                     9762 => "00000001",
                     9763 => "01100110",
                     9764 => "00000000",
                     9765 => "10100111",
                     9766 => "00100010",
                     9767 => "00001000",
                     9768 => "11110010",
                     9769 => "01100111",
                     9770 => "01111011",
                     9771 => "11011100",
                     9772 => "00000010",
                     9773 => "10011000",
                     9774 => "11110010",
                     9775 => "11010111",
                     9776 => "00100000",
                     9777 => "00111001",
                     9778 => "11110001",
                     9779 => "10011111",
                     9780 => "00110011",
                     9781 => "11011100",
                     9782 => "00100111",
                     9783 => "11011100",
                     9784 => "01010111",
                     9785 => "00100011",
                     9786 => "10000011",
                     9787 => "01010111",
                     9788 => "01100011",
                     9789 => "01101100",
                     9790 => "01010001",
                     9791 => "10000111",
                     9792 => "01100011",
                     9793 => "10011001",
                     9794 => "01100001",
                     9795 => "10100011",
                     9796 => "00000110",
                     9797 => "10110011",
                     9798 => "00100001",
                     9799 => "01110111",
                     9800 => "11110011",
                     9801 => "11110011",
                     9802 => "00100001",
                     9803 => "11110111",
                     9804 => "00101010",
                     9805 => "00010011",
                     9806 => "10000001",
                     9807 => "00100011",
                     9808 => "00100010",
                     9809 => "01010011",
                     9810 => "00000000",
                     9811 => "01100011",
                     9812 => "00100010",
                     9813 => "11101001",
                     9814 => "00001011",
                     9815 => "00001100",
                     9816 => "10000011",
                     9817 => "00010011",
                     9818 => "00100001",
                     9819 => "00010110",
                     9820 => "00100010",
                     9821 => "00110011",
                     9822 => "00000101",
                     9823 => "10001111",
                     9824 => "00110101",
                     9825 => "11101100",
                     9826 => "00000001",
                     9827 => "01100011",
                     9828 => "10100000",
                     9829 => "01100111",
                     9830 => "00100000",
                     9831 => "01110011",
                     9832 => "00000001",
                     9833 => "01110111",
                     9834 => "00000001",
                     9835 => "10000011",
                     9836 => "00100000",
                     9837 => "10000111",
                     9838 => "00100000",
                     9839 => "10110011",
                     9840 => "00100000",
                     9841 => "10110111",
                     9842 => "00100000",
                     9843 => "11000011",
                     9844 => "00000001",
                     9845 => "11000111",
                     9846 => "00000000",
                     9847 => "11010011",
                     9848 => "00100000",
                     9849 => "11010111",
                     9850 => "00100000",
                     9851 => "01100111",
                     9852 => "10100000",
                     9853 => "01110111",
                     9854 => "00000111",
                     9855 => "10000111",
                     9856 => "00100010",
                     9857 => "11101000",
                     9858 => "01100010",
                     9859 => "11110101",
                     9860 => "01100101",
                     9861 => "00011100",
                     9862 => "10000010",
                     9863 => "01111111",
                     9864 => "00111000",
                     9865 => "10001101",
                     9866 => "11000001",
                     9867 => "11001111",
                     9868 => "00100110",
                     9869 => "11111101",
                     9870 => "01010000",
                     9871 => "00100001",
                     9872 => "00000111",
                     9873 => "10000001",
                     9874 => "01000111",
                     9875 => "00100100",
                     9876 => "01010111",
                     9877 => "00000000",
                     9878 => "01100011",
                     9879 => "00000001",
                     9880 => "01110111",
                     9881 => "00000001",
                     9882 => "11001001",
                     9883 => "01110001",
                     9884 => "01101000",
                     9885 => "11110010",
                     9886 => "11100111",
                     9887 => "01110011",
                     9888 => "10010111",
                     9889 => "11111011",
                     9890 => "00000110",
                     9891 => "10000011",
                     9892 => "01011100",
                     9893 => "00000001",
                     9894 => "11010111",
                     9895 => "00100010",
                     9896 => "11100111",
                     9897 => "00000000",
                     9898 => "00000011",
                     9899 => "10100111",
                     9900 => "01101100",
                     9901 => "00000010",
                     9902 => "10110011",
                     9903 => "00100010",
                     9904 => "11100011",
                     9905 => "00000001",
                     9906 => "11100111",
                     9907 => "00000111",
                     9908 => "01000111",
                     9909 => "10100000",
                     9910 => "01010111",
                     9911 => "00000110",
                     9912 => "10100111",
                     9913 => "00000001",
                     9914 => "11010011",
                     9915 => "00000000",
                     9916 => "11010111",
                     9917 => "00000001",
                     9918 => "00000111",
                     9919 => "10000001",
                     9920 => "01100111",
                     9921 => "00100000",
                     9922 => "10010011",
                     9923 => "00100010",
                     9924 => "00000011",
                     9925 => "10100011",
                     9926 => "00011100",
                     9927 => "01100001",
                     9928 => "00010111",
                     9929 => "00100001",
                     9930 => "01101111",
                     9931 => "00110011",
                     9932 => "11000111",
                     9933 => "01100011",
                     9934 => "11011000",
                     9935 => "01100010",
                     9936 => "11101001",
                     9937 => "01100001",
                     9938 => "11111010",
                     9939 => "01100000",
                     9940 => "01001111",
                     9941 => "10110011",
                     9942 => "10000111",
                     9943 => "01100011",
                     9944 => "10011100",
                     9945 => "00000001",
                     9946 => "10110111",
                     9947 => "01100011",
                     9948 => "11001000",
                     9949 => "01100010",
                     9950 => "11011001",
                     9951 => "01100001",
                     9952 => "11101010",
                     9953 => "01100000",
                     9954 => "00111001",
                     9955 => "11110001",
                     9956 => "10000111",
                     9957 => "00100001",
                     9958 => "10100111",
                     9959 => "00000001",
                     9960 => "10110111",
                     9961 => "00100000",
                     9962 => "00111001",
                     9963 => "11110001",
                     9964 => "01011111",
                     9965 => "00111000",
                     9966 => "01101101",
                     9967 => "11000001",
                     9968 => "10101111",
                     9969 => "00100110",
                     9970 => "11111101",
                     9971 => "10010000",
                     9972 => "00010001",
                     9973 => "00001111",
                     9974 => "00100110",
                     9975 => "11111110",
                     9976 => "00010000",
                     9977 => "00101010",
                     9978 => "10010011",
                     9979 => "10000111",
                     9980 => "00010111",
                     9981 => "10100011",
                     9982 => "00010100",
                     9983 => "10110010",
                     9984 => "01000010",
                     9985 => "00001010",
                     9986 => "10010010",
                     9987 => "00011001",
                     9988 => "01000000",
                     9989 => "00110110",
                     9990 => "00010100",
                     9991 => "01010000",
                     9992 => "01000001",
                     9993 => "10000010",
                     9994 => "00010110",
                     9995 => "00101011",
                     9996 => "10010011",
                     9997 => "00100100",
                     9998 => "01000001",
                     9999 => "10111011",
                     10000 => "00010100",
                     10001 => "10111000",
                     10002 => "00000000",
                     10003 => "11000010",
                     10004 => "01000011",
                     10005 => "11000011",
                     10006 => "00010011",
                     10007 => "00011011",
                     10008 => "10010100",
                     10009 => "01100111",
                     10010 => "00010010",
                     10011 => "11000100",
                     10012 => "00010101",
                     10013 => "01010011",
                     10014 => "11000001",
                     10015 => "11010010",
                     10016 => "01000001",
                     10017 => "00010010",
                     10018 => "11000001",
                     10019 => "00101001",
                     10020 => "00010011",
                     10021 => "10000101",
                     10022 => "00010111",
                     10023 => "00011011",
                     10024 => "10010010",
                     10025 => "00011010",
                     10026 => "01000010",
                     10027 => "01000111",
                     10028 => "00010011",
                     10029 => "10000011",
                     10030 => "01000001",
                     10031 => "10100111",
                     10032 => "00010011",
                     10033 => "00001110",
                     10034 => "10010001",
                     10035 => "10100111",
                     10036 => "01100011",
                     10037 => "10110111",
                     10038 => "01100011",
                     10039 => "11000101",
                     10040 => "01100101",
                     10041 => "11010101",
                     10042 => "01100101",
                     10043 => "11011101",
                     10044 => "01001010",
                     10045 => "11100011",
                     10046 => "01100111",
                     10047 => "11110011",
                     10048 => "01100111",
                     10049 => "10001101",
                     10050 => "11000001",
                     10051 => "10101110",
                     10052 => "01000010",
                     10053 => "11011111",
                     10054 => "00100000",
                     10055 => "11111101",
                     10056 => "10010000",
                     10057 => "00010001",
                     10058 => "00001111",
                     10059 => "00100110",
                     10060 => "01101110",
                     10061 => "00010000",
                     10062 => "10001011",
                     10063 => "00010111",
                     10064 => "10101111",
                     10065 => "00110010",
                     10066 => "11011000",
                     10067 => "01100010",
                     10068 => "11101000",
                     10069 => "01100010",
                     10070 => "11111100",
                     10071 => "00111111",
                     10072 => "10101101",
                     10073 => "11001000",
                     10074 => "11111000",
                     10075 => "01100100",
                     10076 => "00001100",
                     10077 => "10111110",
                     10078 => "01000011",
                     10079 => "01000011",
                     10080 => "11111000",
                     10081 => "01100100",
                     10082 => "00001100",
                     10083 => "10111111",
                     10084 => "01110011",
                     10085 => "01000000",
                     10086 => "10000100",
                     10087 => "01000000",
                     10088 => "10010011",
                     10089 => "01000000",
                     10090 => "10100100",
                     10091 => "01000000",
                     10092 => "10110011",
                     10093 => "01000000",
                     10094 => "11111000",
                     10095 => "01100100",
                     10096 => "01001000",
                     10097 => "11100100",
                     10098 => "01011100",
                     10099 => "00111001",
                     10100 => "10000011",
                     10101 => "01000000",
                     10102 => "10010010",
                     10103 => "01000001",
                     10104 => "10110011",
                     10105 => "01000000",
                     10106 => "11111000",
                     10107 => "01100100",
                     10108 => "01001000",
                     10109 => "11100100",
                     10110 => "01011100",
                     10111 => "00111001",
                     10112 => "11111000",
                     10113 => "01100100",
                     10114 => "00010011",
                     10115 => "11000010",
                     10116 => "00110111",
                     10117 => "01100101",
                     10118 => "01001100",
                     10119 => "00100100",
                     10120 => "01100011",
                     10121 => "00000000",
                     10122 => "10010111",
                     10123 => "01100101",
                     10124 => "11000011",
                     10125 => "01000010",
                     10126 => "00001011",
                     10127 => "10010111",
                     10128 => "10101100",
                     10129 => "00110010",
                     10130 => "11111000",
                     10131 => "01100100",
                     10132 => "00001100",
                     10133 => "10111110",
                     10134 => "01010011",
                     10135 => "01000101",
                     10136 => "10011101",
                     10137 => "01001000",
                     10138 => "11111000",
                     10139 => "01100100",
                     10140 => "00101010",
                     10141 => "11100010",
                     10142 => "00111100",
                     10143 => "01000111",
                     10144 => "01010110",
                     10145 => "01000011",
                     10146 => "10111010",
                     10147 => "01100010",
                     10148 => "11111000",
                     10149 => "01100100",
                     10150 => "00001100",
                     10151 => "10110111",
                     10152 => "10001000",
                     10153 => "01100100",
                     10154 => "10111100",
                     10155 => "00110001",
                     10156 => "11010100",
                     10157 => "01000101",
                     10158 => "11111100",
                     10159 => "00110001",
                     10160 => "00111100",
                     10161 => "10110001",
                     10162 => "01111000",
                     10163 => "01100100",
                     10164 => "10001100",
                     10165 => "00111000",
                     10166 => "00001011",
                     10167 => "10011100",
                     10168 => "00011010",
                     10169 => "00110011",
                     10170 => "00011000",
                     10171 => "01100001",
                     10172 => "00101000",
                     10173 => "01100001",
                     10174 => "00111001",
                     10175 => "01100000",
                     10176 => "01011101",
                     10177 => "01001010",
                     10178 => "11101110",
                     10179 => "00010001",
                     10180 => "00001111",
                     10181 => "10111000",
                     10182 => "00011101",
                     10183 => "11000001",
                     10184 => "00111110",
                     10185 => "01000010",
                     10186 => "01101111",
                     10187 => "00100000",
                     10188 => "11111101",
                     10189 => "01010010",
                     10190 => "00110001",
                     10191 => "00001111",
                     10192 => "00100000",
                     10193 => "01101110",
                     10194 => "01000000",
                     10195 => "11110111",
                     10196 => "00100000",
                     10197 => "00000111",
                     10198 => "10000100",
                     10199 => "00010111",
                     10200 => "00100000",
                     10201 => "01001111",
                     10202 => "00110100",
                     10203 => "11000011",
                     10204 => "00000011",
                     10205 => "11000111",
                     10206 => "00000010",
                     10207 => "11010011",
                     10208 => "00100010",
                     10209 => "00100111",
                     10210 => "11100011",
                     10211 => "00111001",
                     10212 => "01100001",
                     10213 => "11100111",
                     10214 => "01110011",
                     10215 => "01011100",
                     10216 => "11100100",
                     10217 => "01010111",
                     10218 => "00000000",
                     10219 => "01101100",
                     10220 => "01110011",
                     10221 => "01000111",
                     10222 => "10100000",
                     10223 => "01010011",
                     10224 => "00000110",
                     10225 => "01100011",
                     10226 => "00100010",
                     10227 => "10100111",
                     10228 => "01110011",
                     10229 => "11111100",
                     10230 => "01110011",
                     10231 => "00010011",
                     10232 => "10100001",
                     10233 => "00110011",
                     10234 => "00000101",
                     10235 => "01000011",
                     10236 => "00100001",
                     10237 => "01011100",
                     10238 => "01110010",
                     10239 => "11000011",
                     10240 => "00100011",
                     10241 => "11001100",
                     10242 => "00000011",
                     10243 => "01110111",
                     10244 => "11111011",
                     10245 => "10101100",
                     10246 => "00000010",
                     10247 => "00111001",
                     10248 => "11110001",
                     10249 => "10100111",
                     10250 => "01110011",
                     10251 => "11010011",
                     10252 => "00000100",
                     10253 => "11101000",
                     10254 => "01110010",
                     10255 => "11100011",
                     10256 => "00100010",
                     10257 => "00100110",
                     10258 => "11110100",
                     10259 => "10111100",
                     10260 => "00000010",
                     10261 => "10001100",
                     10262 => "10000001",
                     10263 => "10101000",
                     10264 => "01100010",
                     10265 => "00010111",
                     10266 => "10000111",
                     10267 => "01000011",
                     10268 => "00100100",
                     10269 => "10100111",
                     10270 => "00000001",
                     10271 => "11000011",
                     10272 => "00000100",
                     10273 => "00001000",
                     10274 => "11110010",
                     10275 => "10010111",
                     10276 => "00100001",
                     10277 => "10100011",
                     10278 => "00000010",
                     10279 => "11001001",
                     10280 => "00001011",
                     10281 => "11100001",
                     10282 => "01101001",
                     10283 => "11110001",
                     10284 => "01101001",
                     10285 => "10001101",
                     10286 => "11000001",
                     10287 => "11001111",
                     10288 => "00100110",
                     10289 => "11111101",
                     10290 => "00111000",
                     10291 => "00010001",
                     10292 => "00001111",
                     10293 => "00100110",
                     10294 => "10101101",
                     10295 => "01000000",
                     10296 => "00111101",
                     10297 => "11000111",
                     10298 => "11111101",
                     10299 => "10010101",
                     10300 => "10110001",
                     10301 => "00001111",
                     10302 => "00100110",
                     10303 => "00001101",
                     10304 => "00000010",
                     10305 => "11001000",
                     10306 => "01110010",
                     10307 => "00011100",
                     10308 => "10000001",
                     10309 => "00111000",
                     10310 => "01110010",
                     10311 => "00001101",
                     10312 => "00000101",
                     10313 => "10010111",
                     10314 => "00110100",
                     10315 => "10011000",
                     10316 => "01100010",
                     10317 => "10100011",
                     10318 => "00100000",
                     10319 => "10110011",
                     10320 => "00000110",
                     10321 => "11000011",
                     10322 => "00100000",
                     10323 => "11001100",
                     10324 => "00000011",
                     10325 => "11111001",
                     10326 => "10010001",
                     10327 => "00101100",
                     10328 => "10000001",
                     10329 => "01001000",
                     10330 => "01100010",
                     10331 => "00001101",
                     10332 => "00001001",
                     10333 => "00110111",
                     10334 => "01100011",
                     10335 => "01000111",
                     10336 => "00000011",
                     10337 => "01010111",
                     10338 => "00100001",
                     10339 => "10001100",
                     10340 => "00000010",
                     10341 => "11000101",
                     10342 => "01111001",
                     10343 => "11000111",
                     10344 => "00110001",
                     10345 => "11111001",
                     10346 => "00010001",
                     10347 => "00111001",
                     10348 => "11110001",
                     10349 => "10101001",
                     10350 => "00010001",
                     10351 => "01101111",
                     10352 => "10110100",
                     10353 => "11010011",
                     10354 => "01100101",
                     10355 => "11100011",
                     10356 => "01100101",
                     10357 => "01111101",
                     10358 => "11000001",
                     10359 => "10111111",
                     10360 => "00100110",
                     10361 => "11111101",
                     10362 => "00000000",
                     10363 => "11000001",
                     10364 => "01001100",
                     10365 => "00000000",
                     10366 => "11110100",
                     10367 => "01001111",
                     10368 => "00001101",
                     10369 => "00000010",
                     10370 => "00000010",
                     10371 => "01000010",
                     10372 => "01000011",
                     10373 => "01001111",
                     10374 => "01010010",
                     10375 => "11000010",
                     10376 => "11011110",
                     10377 => "00000000",
                     10378 => "01011010",
                     10379 => "11000010",
                     10380 => "01001101",
                     10381 => "11000111",
                     10382 => "11111101",
                     10383 => "10010000",
                     10384 => "01010001",
                     10385 => "00001111",
                     10386 => "00100110",
                     10387 => "11101110",
                     10388 => "00010000",
                     10389 => "00001011",
                     10390 => "10010100",
                     10391 => "00110011",
                     10392 => "00010100",
                     10393 => "01000010",
                     10394 => "01000010",
                     10395 => "01110111",
                     10396 => "00010110",
                     10397 => "10000110",
                     10398 => "01000100",
                     10399 => "00000010",
                     10400 => "10010010",
                     10401 => "01001010",
                     10402 => "00010110",
                     10403 => "01101001",
                     10404 => "01000010",
                     10405 => "01110011",
                     10406 => "00010100",
                     10407 => "10110000",
                     10408 => "00000000",
                     10409 => "11000111",
                     10410 => "00010010",
                     10411 => "00000101",
                     10412 => "11000000",
                     10413 => "00011100",
                     10414 => "00010111",
                     10415 => "00011111",
                     10416 => "00010001",
                     10417 => "00110110",
                     10418 => "00010010",
                     10419 => "10001111",
                     10420 => "00010100",
                     10421 => "10010001",
                     10422 => "01000000",
                     10423 => "00011011",
                     10424 => "10010100",
                     10425 => "00110101",
                     10426 => "00010010",
                     10427 => "00110100",
                     10428 => "01000010",
                     10429 => "01100000",
                     10430 => "01000010",
                     10431 => "01100001",
                     10432 => "00010010",
                     10433 => "10000111",
                     10434 => "00010010",
                     10435 => "10010110",
                     10436 => "01000000",
                     10437 => "10100011",
                     10438 => "00010100",
                     10439 => "00011100",
                     10440 => "10011000",
                     10441 => "00011111",
                     10442 => "00010001",
                     10443 => "01000111",
                     10444 => "00010010",
                     10445 => "10011111",
                     10446 => "00010101",
                     10447 => "11001100",
                     10448 => "00010101",
                     10449 => "11001111",
                     10450 => "00010001",
                     10451 => "00000101",
                     10452 => "11000000",
                     10453 => "00011111",
                     10454 => "00010101",
                     10455 => "00111001",
                     10456 => "00010010",
                     10457 => "01111100",
                     10458 => "00010110",
                     10459 => "01111111",
                     10460 => "00010001",
                     10461 => "10000010",
                     10462 => "01000000",
                     10463 => "10011000",
                     10464 => "00010010",
                     10465 => "11011111",
                     10466 => "00010101",
                     10467 => "00010110",
                     10468 => "11000100",
                     10469 => "00010111",
                     10470 => "00010100",
                     10471 => "01010100",
                     10472 => "00010010",
                     10473 => "10011011",
                     10474 => "00010110",
                     10475 => "00101000",
                     10476 => "10010100",
                     10477 => "11001110",
                     10478 => "00000001",
                     10479 => "00111101",
                     10480 => "11000001",
                     10481 => "01011110",
                     10482 => "01000010",
                     10483 => "10001111",
                     10484 => "00100000",
                     10485 => "11111101",
                     10486 => "10010111",
                     10487 => "00010001",
                     10488 => "00001111",
                     10489 => "00100110",
                     10490 => "11111110",
                     10491 => "00010000",
                     10492 => "00101011",
                     10493 => "10010010",
                     10494 => "01010111",
                     10495 => "00010010",
                     10496 => "10001011",
                     10497 => "00010010",
                     10498 => "11000000",
                     10499 => "01000001",
                     10500 => "11110111",
                     10501 => "00010011",
                     10502 => "01011011",
                     10503 => "10010010",
                     10504 => "01101001",
                     10505 => "00001011",
                     10506 => "10111011",
                     10507 => "00010010",
                     10508 => "10110010",
                     10509 => "01000110",
                     10510 => "00011001",
                     10511 => "10010011",
                     10512 => "01110001",
                     10513 => "00000000",
                     10514 => "00010111",
                     10515 => "10010100",
                     10516 => "01111100",
                     10517 => "00010100",
                     10518 => "01111111",
                     10519 => "00010001",
                     10520 => "10010011",
                     10521 => "01000001",
                     10522 => "10111111",
                     10523 => "00010101",
                     10524 => "11111100",
                     10525 => "00010011",
                     10526 => "11111111",
                     10527 => "00010001",
                     10528 => "00101111",
                     10529 => "10010101",
                     10530 => "01010000",
                     10531 => "01000010",
                     10532 => "01010001",
                     10533 => "00010010",
                     10534 => "01011000",
                     10535 => "00010100",
                     10536 => "10100110",
                     10537 => "00010010",
                     10538 => "11011011",
                     10539 => "00010010",
                     10540 => "00011011",
                     10541 => "10010011",
                     10542 => "01000110",
                     10543 => "01000011",
                     10544 => "01111011",
                     10545 => "00010010",
                     10546 => "10001101",
                     10547 => "01001001",
                     10548 => "10110111",
                     10549 => "00010100",
                     10550 => "00011011",
                     10551 => "10010100",
                     10552 => "01001001",
                     10553 => "00001011",
                     10554 => "10111011",
                     10555 => "00010010",
                     10556 => "11111100",
                     10557 => "00010011",
                     10558 => "11111111",
                     10559 => "00010010",
                     10560 => "00000011",
                     10561 => "11000001",
                     10562 => "00101111",
                     10563 => "00010101",
                     10564 => "01000011",
                     10565 => "00010010",
                     10566 => "01001011",
                     10567 => "00010011",
                     10568 => "01110111",
                     10569 => "00010011",
                     10570 => "10011101",
                     10571 => "01001010",
                     10572 => "00010101",
                     10573 => "11000001",
                     10574 => "10100001",
                     10575 => "01000001",
                     10576 => "11000011",
                     10577 => "00010010",
                     10578 => "11111110",
                     10579 => "00000001",
                     10580 => "01111101",
                     10581 => "11000001",
                     10582 => "10011110",
                     10583 => "01000010",
                     10584 => "11001111",
                     10585 => "00100000",
                     10586 => "11111101",
                     10587 => "01010010",
                     10588 => "00100001",
                     10589 => "00001111",
                     10590 => "00100000",
                     10591 => "01101110",
                     10592 => "01000100",
                     10593 => "00001100",
                     10594 => "11110001",
                     10595 => "01001100",
                     10596 => "00000001",
                     10597 => "10101010",
                     10598 => "00110101",
                     10599 => "11011001",
                     10600 => "00110100",
                     10601 => "11101110",
                     10602 => "00100000",
                     10603 => "00001000",
                     10604 => "10110011",
                     10605 => "00110111",
                     10606 => "00110010",
                     10607 => "01000011",
                     10608 => "00000100",
                     10609 => "01001110",
                     10610 => "00100001",
                     10611 => "01010011",
                     10612 => "00100000",
                     10613 => "01111100",
                     10614 => "00000001",
                     10615 => "10010111",
                     10616 => "00100001",
                     10617 => "10110111",
                     10618 => "00000111",
                     10619 => "10011100",
                     10620 => "10000001",
                     10621 => "11100111",
                     10622 => "01000010",
                     10623 => "01011111",
                     10624 => "10110011",
                     10625 => "10010111",
                     10626 => "01100011",
                     10627 => "10101100",
                     10628 => "00000010",
                     10629 => "11000101",
                     10630 => "01000001",
                     10631 => "01001001",
                     10632 => "11100000",
                     10633 => "01011000",
                     10634 => "01100001",
                     10635 => "01110110",
                     10636 => "01100100",
                     10637 => "10000101",
                     10638 => "01100101",
                     10639 => "10010100",
                     10640 => "01100110",
                     10641 => "10100100",
                     10642 => "00100010",
                     10643 => "10100110",
                     10644 => "00000011",
                     10645 => "11001000",
                     10646 => "00100010",
                     10647 => "11011100",
                     10648 => "00000010",
                     10649 => "01101000",
                     10650 => "11110010",
                     10651 => "10010110",
                     10652 => "01000010",
                     10653 => "00010011",
                     10654 => "10000010",
                     10655 => "00010111",
                     10656 => "00000010",
                     10657 => "10101111",
                     10658 => "00110100",
                     10659 => "11110110",
                     10660 => "00100001",
                     10661 => "11111100",
                     10662 => "00000110",
                     10663 => "00100110",
                     10664 => "10000000",
                     10665 => "00101010",
                     10666 => "00100100",
                     10667 => "00110110",
                     10668 => "00000001",
                     10669 => "10001100",
                     10670 => "00000000",
                     10671 => "11111111",
                     10672 => "00110101",
                     10673 => "01001110",
                     10674 => "10100000",
                     10675 => "01010101",
                     10676 => "00100001",
                     10677 => "01110111",
                     10678 => "00100000",
                     10679 => "10000111",
                     10680 => "00000111",
                     10681 => "10001001",
                     10682 => "00100010",
                     10683 => "10101110",
                     10684 => "00100001",
                     10685 => "01001100",
                     10686 => "10000010",
                     10687 => "10011111",
                     10688 => "00110100",
                     10689 => "11101100",
                     10690 => "00000001",
                     10691 => "00000011",
                     10692 => "11100111",
                     10693 => "00010011",
                     10694 => "01100111",
                     10695 => "10001101",
                     10696 => "01001010",
                     10697 => "10101101",
                     10698 => "01000001",
                     10699 => "00001111",
                     10700 => "10100110",
                     10701 => "11111101",
                     10702 => "00010000",
                     10703 => "01010001",
                     10704 => "01001100",
                     10705 => "00000000",
                     10706 => "11000111",
                     10707 => "00010010",
                     10708 => "11000110",
                     10709 => "01000010",
                     10710 => "00000011",
                     10711 => "10010010",
                     10712 => "00000010",
                     10713 => "01000010",
                     10714 => "00101001",
                     10715 => "00010010",
                     10716 => "01100011",
                     10717 => "00010010",
                     10718 => "01100010",
                     10719 => "01000010",
                     10720 => "01101001",
                     10721 => "00010100",
                     10722 => "10100101",
                     10723 => "00010010",
                     10724 => "10100100",
                     10725 => "01000010",
                     10726 => "11100010",
                     10727 => "00010100",
                     10728 => "11100001",
                     10729 => "01000100",
                     10730 => "11111000",
                     10731 => "00010110",
                     10732 => "00110111",
                     10733 => "11000001",
                     10734 => "10001111",
                     10735 => "00111000",
                     10736 => "00000010",
                     10737 => "10111011",
                     10738 => "00101000",
                     10739 => "01111010",
                     10740 => "01101000",
                     10741 => "01111010",
                     10742 => "10101000",
                     10743 => "01111010",
                     10744 => "11100000",
                     10745 => "01101010",
                     10746 => "11110000",
                     10747 => "01101010",
                     10748 => "01101101",
                     10749 => "11000101",
                     10750 => "11111101",
                     10751 => "10010010",
                     10752 => "00110001",
                     10753 => "00001111",
                     10754 => "00100000",
                     10755 => "01101110",
                     10756 => "01000000",
                     10757 => "00001101",
                     10758 => "00000010",
                     10759 => "00110111",
                     10760 => "01110011",
                     10761 => "11101100",
                     10762 => "00000000",
                     10763 => "00001100",
                     10764 => "10000000",
                     10765 => "00111100",
                     10766 => "00000000",
                     10767 => "01101100",
                     10768 => "00000000",
                     10769 => "10011100",
                     10770 => "00000000",
                     10771 => "00000110",
                     10772 => "11000000",
                     10773 => "11000111",
                     10774 => "01110011",
                     10775 => "00000110",
                     10776 => "10000011",
                     10777 => "00101000",
                     10778 => "01110010",
                     10779 => "10010110",
                     10780 => "01000000",
                     10781 => "11100111",
                     10782 => "01110011",
                     10783 => "00100110",
                     10784 => "11000000",
                     10785 => "10000111",
                     10786 => "01111011",
                     10787 => "11010010",
                     10788 => "01000001",
                     10789 => "00111001",
                     10790 => "11110001",
                     10791 => "11001000",
                     10792 => "11110010",
                     10793 => "10010111",
                     10794 => "11100011",
                     10795 => "10100011",
                     10796 => "00100011",
                     10797 => "11100111",
                     10798 => "00000010",
                     10799 => "11100011",
                     10800 => "00000111",
                     10801 => "11110011",
                     10802 => "00100010",
                     10803 => "00110111",
                     10804 => "11100011",
                     10805 => "10011100",
                     10806 => "00000000",
                     10807 => "10111100",
                     10808 => "00000000",
                     10809 => "11101100",
                     10810 => "00000000",
                     10811 => "00001100",
                     10812 => "10000000",
                     10813 => "00111100",
                     10814 => "00000000",
                     10815 => "10000110",
                     10816 => "00100001",
                     10817 => "10100110",
                     10818 => "00000110",
                     10819 => "10110110",
                     10820 => "00100100",
                     10821 => "01011100",
                     10822 => "10000000",
                     10823 => "01111100",
                     10824 => "00000000",
                     10825 => "10011100",
                     10826 => "00000000",
                     10827 => "00101001",
                     10828 => "11100001",
                     10829 => "11011100",
                     10830 => "00000101",
                     10831 => "11110110",
                     10832 => "01000001",
                     10833 => "11011100",
                     10834 => "10000000",
                     10835 => "11101000",
                     10836 => "01110010",
                     10837 => "00001100",
                     10838 => "10000001",
                     10839 => "00100111",
                     10840 => "01110011",
                     10841 => "01001100",
                     10842 => "00000001",
                     10843 => "01100110",
                     10844 => "01110100",
                     10845 => "00001101",
                     10846 => "00010001",
                     10847 => "00111111",
                     10848 => "00110101",
                     10849 => "10110110",
                     10850 => "01000001",
                     10851 => "00101100",
                     10852 => "10000010",
                     10853 => "00110110",
                     10854 => "01000000",
                     10855 => "01111100",
                     10856 => "00000010",
                     10857 => "10000110",
                     10858 => "01000000",
                     10859 => "11111001",
                     10860 => "01100001",
                     10861 => "00111001",
                     10862 => "11100001",
                     10863 => "10101100",
                     10864 => "00000100",
                     10865 => "11000110",
                     10866 => "01000001",
                     10867 => "00001100",
                     10868 => "10000011",
                     10869 => "00010110",
                     10870 => "01000001",
                     10871 => "10001000",
                     10872 => "11110010",
                     10873 => "00111001",
                     10874 => "11110001",
                     10875 => "01111100",
                     10876 => "00000000",
                     10877 => "10001001",
                     10878 => "01100001",
                     10879 => "10011100",
                     10880 => "00000000",
                     10881 => "10100111",
                     10882 => "01100011",
                     10883 => "10111100",
                     10884 => "00000000",
                     10885 => "11000101",
                     10886 => "01100101",
                     10887 => "11011100",
                     10888 => "00000000",
                     10889 => "11100011",
                     10890 => "01100111",
                     10891 => "11110011",
                     10892 => "01100111",
                     10893 => "10001101",
                     10894 => "11000001",
                     10895 => "11001111",
                     10896 => "00100110",
                     10897 => "11111101",
                     10898 => "01010101",
                     10899 => "10110001",
                     10900 => "00001111",
                     10901 => "00100110",
                     10902 => "11001111",
                     10903 => "00110011",
                     10904 => "00000111",
                     10905 => "10110010",
                     10906 => "00010101",
                     10907 => "00010001",
                     10908 => "01010010",
                     10909 => "01000010",
                     10910 => "10011001",
                     10911 => "00001011",
                     10912 => "10101100",
                     10913 => "00000010",
                     10914 => "11010011",
                     10915 => "00100100",
                     10916 => "11010110",
                     10917 => "01000010",
                     10918 => "11010111",
                     10919 => "00100101",
                     10920 => "00100011",
                     10921 => "10000100",
                     10922 => "11001111",
                     10923 => "00110011",
                     10924 => "00000111",
                     10925 => "11100011",
                     10926 => "00011001",
                     10927 => "01100001",
                     10928 => "01111000",
                     10929 => "01111010",
                     10930 => "11101111",
                     10931 => "00110011",
                     10932 => "00101100",
                     10933 => "10000001",
                     10934 => "01000110",
                     10935 => "01100100",
                     10936 => "01010101",
                     10937 => "01100101",
                     10938 => "01100101",
                     10939 => "01100101",
                     10940 => "11101100",
                     10941 => "01110100",
                     10942 => "01000111",
                     10943 => "10000010",
                     10944 => "01010011",
                     10945 => "00000101",
                     10946 => "01100011",
                     10947 => "00100001",
                     10948 => "01100010",
                     10949 => "01000001",
                     10950 => "10010110",
                     10951 => "00100010",
                     10952 => "10011010",
                     10953 => "01000001",
                     10954 => "11001100",
                     10955 => "00000011",
                     10956 => "10111001",
                     10957 => "10010001",
                     10958 => "00111001",
                     10959 => "11110001",
                     10960 => "01100011",
                     10961 => "00100110",
                     10962 => "01100111",
                     10963 => "00100111",
                     10964 => "11010011",
                     10965 => "00000110",
                     10966 => "11111100",
                     10967 => "00000001",
                     10968 => "00011000",
                     10969 => "11100010",
                     10970 => "11011001",
                     10971 => "00000111",
                     10972 => "11101001",
                     10973 => "00000100",
                     10974 => "00001100",
                     10975 => "10000110",
                     10976 => "00110111",
                     10977 => "00100010",
                     10978 => "10010011",
                     10979 => "00100100",
                     10980 => "10000111",
                     10981 => "10000100",
                     10982 => "10101100",
                     10983 => "00000010",
                     10984 => "11000010",
                     10985 => "01000001",
                     10986 => "11000011",
                     10987 => "00100011",
                     10988 => "11011001",
                     10989 => "01110001",
                     10990 => "11111100",
                     10991 => "00000001",
                     10992 => "01111111",
                     10993 => "10110001",
                     10994 => "10011100",
                     10995 => "00000000",
                     10996 => "10100111",
                     10997 => "01100011",
                     10998 => "10110110",
                     10999 => "01100100",
                     11000 => "11001100",
                     11001 => "00000000",
                     11002 => "11010100",
                     11003 => "01100110",
                     11004 => "11100011",
                     11005 => "01100111",
                     11006 => "11110011",
                     11007 => "01100111",
                     11008 => "10001101",
                     11009 => "11000001",
                     11010 => "11001111",
                     11011 => "00100110",
                     11012 => "11111101",
                     11013 => "01010000",
                     11014 => "10110001",
                     11015 => "00001111",
                     11016 => "00100110",
                     11017 => "11111100",
                     11018 => "00000000",
                     11019 => "00011111",
                     11020 => "10110011",
                     11021 => "01011100",
                     11022 => "00000000",
                     11023 => "01100101",
                     11024 => "01100101",
                     11025 => "01110100",
                     11026 => "01100110",
                     11027 => "10000011",
                     11028 => "01100111",
                     11029 => "10010011",
                     11030 => "01100111",
                     11031 => "11011100",
                     11032 => "01110011",
                     11033 => "01001100",
                     11034 => "10000000",
                     11035 => "10110011",
                     11036 => "00100000",
                     11037 => "11001001",
                     11038 => "00001011",
                     11039 => "11000011",
                     11040 => "00001000",
                     11041 => "11010011",
                     11042 => "00101111",
                     11043 => "11011100",
                     11044 => "00000000",
                     11045 => "00101100",
                     11046 => "10000000",
                     11047 => "01001100",
                     11048 => "00000000",
                     11049 => "10001100",
                     11050 => "00000000",
                     11051 => "11010011",
                     11052 => "00101110",
                     11053 => "11101101",
                     11054 => "01001010",
                     11055 => "11111100",
                     11056 => "00000000",
                     11057 => "11010111",
                     11058 => "10100001",
                     11059 => "11101100",
                     11060 => "00000001",
                     11061 => "01001100",
                     11062 => "10000000",
                     11063 => "01011001",
                     11064 => "00010001",
                     11065 => "11011000",
                     11066 => "00010001",
                     11067 => "11011010",
                     11068 => "00010000",
                     11069 => "00110111",
                     11070 => "10100000",
                     11071 => "01000111",
                     11072 => "00000100",
                     11073 => "10011001",
                     11074 => "00010001",
                     11075 => "11100111",
                     11076 => "00100001",
                     11077 => "00111010",
                     11078 => "10010000",
                     11079 => "01100111",
                     11080 => "00100000",
                     11081 => "01110110",
                     11082 => "00010000",
                     11083 => "01110111",
                     11084 => "01100000",
                     11085 => "10000111",
                     11086 => "00000111",
                     11087 => "11011000",
                     11088 => "00010010",
                     11089 => "00111001",
                     11090 => "11110001",
                     11091 => "10101100",
                     11092 => "00000000",
                     11093 => "11101001",
                     11094 => "01110001",
                     11095 => "00001100",
                     11096 => "10000000",
                     11097 => "00101100",
                     11098 => "00000000",
                     11099 => "01001100",
                     11100 => "00000101",
                     11101 => "11000111",
                     11102 => "01111011",
                     11103 => "00111001",
                     11104 => "11110001",
                     11105 => "11101100",
                     11106 => "00000000",
                     11107 => "11111001",
                     11108 => "00010001",
                     11109 => "00001100",
                     11110 => "10000010",
                     11111 => "01101111",
                     11112 => "00110100",
                     11113 => "11111000",
                     11114 => "00010001",
                     11115 => "11111010",
                     11116 => "00010000",
                     11117 => "01111111",
                     11118 => "10110010",
                     11119 => "10101100",
                     11120 => "00000000",
                     11121 => "10110110",
                     11122 => "01100100",
                     11123 => "11001100",
                     11124 => "00000001",
                     11125 => "11100011",
                     11126 => "01100111",
                     11127 => "11110011",
                     11128 => "01100111",
                     11129 => "10001101",
                     11130 => "11000001",
                     11131 => "11001111",
                     11132 => "00100110",
                     11133 => "11111101",
                     11134 => "01010010",
                     11135 => "10110001",
                     11136 => "00001111",
                     11137 => "00100000",
                     11138 => "01101110",
                     11139 => "01000101",
                     11140 => "00111001",
                     11141 => "10010001",
                     11142 => "10110011",
                     11143 => "00000100",
                     11144 => "11000011",
                     11145 => "00100001",
                     11146 => "11001000",
                     11147 => "00010001",
                     11148 => "11001010",
                     11149 => "00010000",
                     11150 => "01001001",
                     11151 => "10010001",
                     11152 => "01111100",
                     11153 => "01110011",
                     11154 => "11101000",
                     11155 => "00010010",
                     11156 => "10001000",
                     11157 => "10010001",
                     11158 => "10001010",
                     11159 => "00010000",
                     11160 => "11100111",
                     11161 => "00100001",
                     11162 => "00000101",
                     11163 => "10010001",
                     11164 => "00000111",
                     11165 => "00110000",
                     11166 => "00010111",
                     11167 => "00000111",
                     11168 => "00100111",
                     11169 => "00100000",
                     11170 => "01001001",
                     11171 => "00010001",
                     11172 => "10011100",
                     11173 => "00000001",
                     11174 => "11001000",
                     11175 => "01110010",
                     11176 => "00100011",
                     11177 => "10100110",
                     11178 => "00100111",
                     11179 => "00100110",
                     11180 => "11010011",
                     11181 => "00000011",
                     11182 => "11011000",
                     11183 => "01111010",
                     11184 => "10001001",
                     11185 => "10010001",
                     11186 => "11011000",
                     11187 => "01110010",
                     11188 => "00111001",
                     11189 => "11110001",
                     11190 => "10101001",
                     11191 => "00010001",
                     11192 => "00001001",
                     11193 => "11110001",
                     11194 => "01100011",
                     11195 => "00100100",
                     11196 => "01100111",
                     11197 => "00100100",
                     11198 => "11011000",
                     11199 => "01100010",
                     11200 => "00101000",
                     11201 => "10010001",
                     11202 => "00101010",
                     11203 => "00010000",
                     11204 => "01010110",
                     11205 => "00100001",
                     11206 => "01110000",
                     11207 => "00000100",
                     11208 => "01111001",
                     11209 => "00001011",
                     11210 => "10001100",
                     11211 => "00000000",
                     11212 => "10010100",
                     11213 => "00100001",
                     11214 => "10011111",
                     11215 => "00110101",
                     11216 => "00101111",
                     11217 => "10111000",
                     11218 => "00111101",
                     11219 => "11000001",
                     11220 => "01111111",
                     11221 => "00100110",
                     11222 => "11111101",
                     11223 => "00000110",
                     11224 => "11000001",
                     11225 => "01001100",
                     11226 => "00000000",
                     11227 => "11110100",
                     11228 => "01001111",
                     11229 => "00001101",
                     11230 => "00000010",
                     11231 => "00000110",
                     11232 => "00100000",
                     11233 => "00100100",
                     11234 => "01001111",
                     11235 => "00110101",
                     11236 => "10100000",
                     11237 => "00110110",
                     11238 => "00100000",
                     11239 => "01010011",
                     11240 => "01000110",
                     11241 => "11010101",
                     11242 => "00100000",
                     11243 => "11010110",
                     11244 => "00100000",
                     11245 => "00110100",
                     11246 => "10100001",
                     11247 => "01110011",
                     11248 => "01001001",
                     11249 => "01110100",
                     11250 => "00100000",
                     11251 => "10010100",
                     11252 => "00100000",
                     11253 => "10110100",
                     11254 => "00100000",
                     11255 => "11010100",
                     11256 => "00100000",
                     11257 => "11110100",
                     11258 => "00100000",
                     11259 => "00101110",
                     11260 => "10000000",
                     11261 => "01011001",
                     11262 => "01000010",
                     11263 => "01001101",
                     11264 => "11000111",
                     11265 => "11111101",
                     11266 => "10010110",
                     11267 => "00110001",
                     11268 => "00001111",
                     11269 => "00100110",
                     11270 => "00001101",
                     11271 => "00000011",
                     11272 => "00011010",
                     11273 => "01100000",
                     11274 => "01110111",
                     11275 => "01000010",
                     11276 => "11000100",
                     11277 => "00000000",
                     11278 => "11001000",
                     11279 => "01100010",
                     11280 => "10111001",
                     11281 => "11100001",
                     11282 => "11010011",
                     11283 => "00000110",
                     11284 => "11010111",
                     11285 => "00000111",
                     11286 => "11111001",
                     11287 => "01100001",
                     11288 => "00001100",
                     11289 => "10000001",
                     11290 => "01001110",
                     11291 => "10110001",
                     11292 => "10001110",
                     11293 => "10110001",
                     11294 => "10111100",
                     11295 => "00000001",
                     11296 => "11100100",
                     11297 => "01010000",
                     11298 => "11101001",
                     11299 => "01100001",
                     11300 => "00001100",
                     11301 => "10000001",
                     11302 => "00001101",
                     11303 => "00001010",
                     11304 => "10000100",
                     11305 => "01000011",
                     11306 => "10011000",
                     11307 => "01110010",
                     11308 => "00001101",
                     11309 => "00001100",
                     11310 => "00001111",
                     11311 => "00111000",
                     11312 => "00011101",
                     11313 => "11000001",
                     11314 => "01011111",
                     11315 => "00100110",
                     11316 => "11111101",
                     11317 => "01001000",
                     11318 => "00001111",
                     11319 => "00001110",
                     11320 => "00000001",
                     11321 => "01011110",
                     11322 => "00000010",
                     11323 => "10100111",
                     11324 => "00000000",
                     11325 => "10111100",
                     11326 => "01110011",
                     11327 => "00011010",
                     11328 => "11100000",
                     11329 => "00111001",
                     11330 => "01100001",
                     11331 => "01011000",
                     11332 => "01100010",
                     11333 => "01110111",
                     11334 => "01100011",
                     11335 => "10010111",
                     11336 => "01100011",
                     11337 => "10111000",
                     11338 => "01100010",
                     11339 => "11010110",
                     11340 => "00000111",
                     11341 => "11111000",
                     11342 => "01100010",
                     11343 => "00011001",
                     11344 => "11100001",
                     11345 => "01110101",
                     11346 => "01010010",
                     11347 => "10000110",
                     11348 => "01000000",
                     11349 => "10000111",
                     11350 => "01010000",
                     11351 => "10010101",
                     11352 => "01010010",
                     11353 => "10010011",
                     11354 => "01000011",
                     11355 => "10100101",
                     11356 => "00100001",
                     11357 => "11000101",
                     11358 => "01010010",
                     11359 => "11010110",
                     11360 => "01000000",
                     11361 => "11010111",
                     11362 => "00100000",
                     11363 => "11100101",
                     11364 => "00000110",
                     11365 => "11100110",
                     11366 => "01010001",
                     11367 => "00111110",
                     11368 => "10001101",
                     11369 => "01011110",
                     11370 => "00000011",
                     11371 => "01100111",
                     11372 => "01010010",
                     11373 => "01110111",
                     11374 => "01010010",
                     11375 => "01111110",
                     11376 => "00000010",
                     11377 => "10011110",
                     11378 => "00000011",
                     11379 => "10100110",
                     11380 => "01000011",
                     11381 => "10100111",
                     11382 => "00100011",
                     11383 => "11011110",
                     11384 => "00000101",
                     11385 => "11111110",
                     11386 => "00000010",
                     11387 => "00011110",
                     11388 => "10000011",
                     11389 => "00110011",
                     11390 => "01010100",
                     11391 => "01000110",
                     11392 => "01000000",
                     11393 => "01000111",
                     11394 => "00100001",
                     11395 => "01010110",
                     11396 => "00000100",
                     11397 => "01011110",
                     11398 => "00000010",
                     11399 => "10000011",
                     11400 => "01010100",
                     11401 => "10010011",
                     11402 => "01010010",
                     11403 => "10010110",
                     11404 => "00000111",
                     11405 => "10010111",
                     11406 => "01010000",
                     11407 => "10111110",
                     11408 => "00000011",
                     11409 => "11000111",
                     11410 => "00100011",
                     11411 => "11111110",
                     11412 => "00000010",
                     11413 => "00001100",
                     11414 => "10000010",
                     11415 => "01000011",
                     11416 => "01000101",
                     11417 => "01000101",
                     11418 => "00100100",
                     11419 => "01000110",
                     11420 => "00100100",
                     11421 => "10010000",
                     11422 => "00001000",
                     11423 => "10010101",
                     11424 => "01010001",
                     11425 => "01111000",
                     11426 => "11111010",
                     11427 => "11010111",
                     11428 => "01110011",
                     11429 => "00111001",
                     11430 => "11110001",
                     11431 => "10001100",
                     11432 => "00000001",
                     11433 => "10101000",
                     11434 => "01010010",
                     11435 => "10111000",
                     11436 => "01010010",
                     11437 => "11001100",
                     11438 => "00000001",
                     11439 => "01011111",
                     11440 => "10110011",
                     11441 => "10010111",
                     11442 => "01100011",
                     11443 => "10011110",
                     11444 => "00000000",
                     11445 => "00001110",
                     11446 => "10000001",
                     11447 => "00010110",
                     11448 => "00100100",
                     11449 => "01100110",
                     11450 => "00000100",
                     11451 => "10001110",
                     11452 => "00000000",
                     11453 => "11111110",
                     11454 => "00000001",
                     11455 => "00001000",
                     11456 => "11010010",
                     11457 => "00001110",
                     11458 => "00000110",
                     11459 => "01101111",
                     11460 => "01000111",
                     11461 => "10011110",
                     11462 => "00001111",
                     11463 => "00001110",
                     11464 => "10000010",
                     11465 => "00101101",
                     11466 => "01000111",
                     11467 => "00101000",
                     11468 => "01111010",
                     11469 => "01101000",
                     11470 => "01111010",
                     11471 => "10101000",
                     11472 => "01111010",
                     11473 => "10101110",
                     11474 => "00000001",
                     11475 => "11011110",
                     11476 => "00001111",
                     11477 => "01101101",
                     11478 => "11000101",
                     11479 => "11111101",
                     11480 => "01001000",
                     11481 => "00001111",
                     11482 => "00001110",
                     11483 => "00000001",
                     11484 => "01011110",
                     11485 => "00000010",
                     11486 => "10111100",
                     11487 => "00000001",
                     11488 => "11111100",
                     11489 => "00000001",
                     11490 => "00101100",
                     11491 => "10000010",
                     11492 => "01000001",
                     11493 => "01010010",
                     11494 => "01001110",
                     11495 => "00000100",
                     11496 => "01100111",
                     11497 => "00100101",
                     11498 => "01101000",
                     11499 => "00100100",
                     11500 => "01101001",
                     11501 => "00100100",
                     11502 => "10111010",
                     11503 => "01000010",
                     11504 => "11000111",
                     11505 => "00000100",
                     11506 => "11011110",
                     11507 => "00001011",
                     11508 => "10110010",
                     11509 => "10000111",
                     11510 => "11111110",
                     11511 => "00000010",
                     11512 => "00101100",
                     11513 => "11100001",
                     11514 => "00101100",
                     11515 => "01110001",
                     11516 => "01100111",
                     11517 => "00000001",
                     11518 => "01110111",
                     11519 => "00000000",
                     11520 => "10000111",
                     11521 => "00000001",
                     11522 => "10001110",
                     11523 => "00000000",
                     11524 => "11101110",
                     11525 => "00000001",
                     11526 => "11110110",
                     11527 => "00000010",
                     11528 => "00000011",
                     11529 => "10000101",
                     11530 => "00000101",
                     11531 => "00000010",
                     11532 => "00010011",
                     11533 => "00100001",
                     11534 => "00010110",
                     11535 => "00000010",
                     11536 => "00100111",
                     11537 => "00000010",
                     11538 => "00101110",
                     11539 => "00000010",
                     11540 => "10001000",
                     11541 => "01110010",
                     11542 => "11000111",
                     11543 => "00100000",
                     11544 => "11010111",
                     11545 => "00000111",
                     11546 => "11100100",
                     11547 => "01110110",
                     11548 => "00000111",
                     11549 => "10100000",
                     11550 => "00010111",
                     11551 => "00000110",
                     11552 => "01001000",
                     11553 => "01111010",
                     11554 => "01110110",
                     11555 => "00100000",
                     11556 => "10011000",
                     11557 => "01110010",
                     11558 => "01111001",
                     11559 => "11100001",
                     11560 => "10001000",
                     11561 => "01100010",
                     11562 => "10011100",
                     11563 => "00000001",
                     11564 => "10110111",
                     11565 => "01110011",
                     11566 => "11011100",
                     11567 => "00000001",
                     11568 => "11111000",
                     11569 => "01100010",
                     11570 => "11111110",
                     11571 => "00000001",
                     11572 => "00001000",
                     11573 => "11100010",
                     11574 => "00001110",
                     11575 => "00000000",
                     11576 => "01101110",
                     11577 => "00000010",
                     11578 => "01110011",
                     11579 => "00100000",
                     11580 => "01110111",
                     11581 => "00100011",
                     11582 => "10000011",
                     11583 => "00000100",
                     11584 => "10010011",
                     11585 => "00100000",
                     11586 => "10101110",
                     11587 => "00000000",
                     11588 => "11111110",
                     11589 => "00001010",
                     11590 => "00001110",
                     11591 => "10000010",
                     11592 => "00111001",
                     11593 => "01110001",
                     11594 => "10101000",
                     11595 => "01110010",
                     11596 => "11100111",
                     11597 => "01110011",
                     11598 => "00001100",
                     11599 => "10000001",
                     11600 => "10001111",
                     11601 => "00110010",
                     11602 => "10101110",
                     11603 => "00000000",
                     11604 => "11111110",
                     11605 => "00000100",
                     11606 => "00000100",
                     11607 => "11010001",
                     11608 => "00010111",
                     11609 => "00000100",
                     11610 => "00100110",
                     11611 => "01001001",
                     11612 => "00100111",
                     11613 => "00101001",
                     11614 => "11011111",
                     11615 => "00110011",
                     11616 => "11111110",
                     11617 => "00000010",
                     11618 => "01000100",
                     11619 => "11110110",
                     11620 => "01111100",
                     11621 => "00000001",
                     11622 => "10001110",
                     11623 => "00000110",
                     11624 => "10111111",
                     11625 => "01000111",
                     11626 => "11101110",
                     11627 => "00001111",
                     11628 => "01001101",
                     11629 => "11000111",
                     11630 => "00001110",
                     11631 => "10000010",
                     11632 => "01101000",
                     11633 => "01111010",
                     11634 => "10101110",
                     11635 => "00000001",
                     11636 => "11011110",
                     11637 => "00001111",
                     11638 => "01101101",
                     11639 => "11000101",
                     11640 => "11111101",
                     11641 => "01001000",
                     11642 => "00000001",
                     11643 => "00001110",
                     11644 => "00000001",
                     11645 => "00000000",
                     11646 => "01011010",
                     11647 => "00111110",
                     11648 => "00000110",
                     11649 => "01000101",
                     11650 => "01000110",
                     11651 => "01000111",
                     11652 => "01000110",
                     11653 => "01010011",
                     11654 => "01000100",
                     11655 => "10101110",
                     11656 => "00000001",
                     11657 => "11011111",
                     11658 => "01001010",
                     11659 => "01001101",
                     11660 => "11000111",
                     11661 => "00001110",
                     11662 => "10000001",
                     11663 => "00000000",
                     11664 => "01011010",
                     11665 => "00101110",
                     11666 => "00000100",
                     11667 => "00110111",
                     11668 => "00101000",
                     11669 => "00111010",
                     11670 => "01001000",
                     11671 => "01000110",
                     11672 => "01000111",
                     11673 => "11000111",
                     11674 => "00000111",
                     11675 => "11001110",
                     11676 => "00001111",
                     11677 => "11011111",
                     11678 => "01001010",
                     11679 => "01001101",
                     11680 => "11000111",
                     11681 => "00001110",
                     11682 => "10000001",
                     11683 => "00000000",
                     11684 => "01011010",
                     11685 => "00110011",
                     11686 => "01010011",
                     11687 => "01000011",
                     11688 => "01010001",
                     11689 => "01000110",
                     11690 => "01000000",
                     11691 => "01000111",
                     11692 => "01010000",
                     11693 => "01010011",
                     11694 => "00000100",
                     11695 => "01010101",
                     11696 => "01000000",
                     11697 => "01010110",
                     11698 => "01010000",
                     11699 => "01100010",
                     11700 => "01000011",
                     11701 => "01100100",
                     11702 => "01000000",
                     11703 => "01100101",
                     11704 => "01010000",
                     11705 => "01110001",
                     11706 => "01000001",
                     11707 => "01110011",
                     11708 => "01010001",
                     11709 => "10000011",
                     11710 => "01010001",
                     11711 => "10010100",
                     11712 => "01000000",
                     11713 => "10010101",
                     11714 => "01010000",
                     11715 => "10100011",
                     11716 => "01010000",
                     11717 => "10100101",
                     11718 => "01000000",
                     11719 => "10100110",
                     11720 => "01010000",
                     11721 => "10110011",
                     11722 => "01010001",
                     11723 => "10110110",
                     11724 => "01000000",
                     11725 => "10110111",
                     11726 => "01010000",
                     11727 => "11000011",
                     11728 => "01010011",
                     11729 => "11011111",
                     11730 => "01001010",
                     11731 => "01001101",
                     11732 => "11000111",
                     11733 => "00001110",
                     11734 => "10000001",
                     11735 => "00000000",
                     11736 => "01011010",
                     11737 => "00101110",
                     11738 => "00000010",
                     11739 => "00110110",
                     11740 => "01000111",
                     11741 => "00110111",
                     11742 => "01010010",
                     11743 => "00111010",
                     11744 => "01001001",
                     11745 => "01000111",
                     11746 => "00100101",
                     11747 => "10100111",
                     11748 => "01010010",
                     11749 => "11010111",
                     11750 => "00000100",
                     11751 => "11011111",
                     11752 => "01001010",
                     11753 => "01001101",
                     11754 => "11000111",
                     11755 => "00001110",
                     11756 => "10000001",
                     11757 => "00000000",
                     11758 => "01011010",
                     11759 => "00111110",
                     11760 => "00000010",
                     11761 => "01000100",
                     11762 => "01010001",
                     11763 => "01010011",
                     11764 => "01000100",
                     11765 => "01010100",
                     11766 => "01000100",
                     11767 => "01010101",
                     11768 => "00100100",
                     11769 => "10100001",
                     11770 => "01010100",
                     11771 => "10101110",
                     11772 => "00000001",
                     11773 => "10110100",
                     11774 => "00100001",
                     11775 => "11011111",
                     11776 => "01001010",
                     11777 => "11100101",
                     11778 => "00000111",
                     11779 => "01001101",
                     11780 => "11000111",
                     11781 => "11111101",
                     11782 => "01000001",
                     11783 => "00000001",
                     11784 => "10110100",
                     11785 => "00110100",
                     11786 => "11001000",
                     11787 => "01010010",
                     11788 => "11110010",
                     11789 => "01010001",
                     11790 => "01000111",
                     11791 => "11010011",
                     11792 => "01101100",
                     11793 => "00000011",
                     11794 => "01100101",
                     11795 => "01001001",
                     11796 => "10011110",
                     11797 => "00000111",
                     11798 => "10111110",
                     11799 => "00000001",
                     11800 => "11001100",
                     11801 => "00000011",
                     11802 => "11111110",
                     11803 => "00000111",
                     11804 => "00001101",
                     11805 => "11001001",
                     11806 => "00011110",
                     11807 => "00000001",
                     11808 => "01101100",
                     11809 => "00000001",
                     11810 => "01100010",
                     11811 => "00110101",
                     11812 => "01100011",
                     11813 => "01010011",
                     11814 => "10001010",
                     11815 => "01000001",
                     11816 => "10101100",
                     11817 => "00000001",
                     11818 => "10110011",
                     11819 => "01010011",
                     11820 => "11101001",
                     11821 => "01010001",
                     11822 => "00100110",
                     11823 => "11000011",
                     11824 => "00100111",
                     11825 => "00110011",
                     11826 => "01100011",
                     11827 => "01000011",
                     11828 => "01100100",
                     11829 => "00110011",
                     11830 => "10111010",
                     11831 => "01100000",
                     11832 => "11001001",
                     11833 => "01100001",
                     11834 => "11001110",
                     11835 => "00001011",
                     11836 => "11011110",
                     11837 => "00001111",
                     11838 => "11100101",
                     11839 => "00001001",
                     11840 => "01111101",
                     11841 => "11001010",
                     11842 => "01111101",
                     11843 => "01000111",
                     11844 => "11111101",
                     11845 => "01000001",
                     11846 => "00000001",
                     11847 => "10111000",
                     11848 => "01010010",
                     11849 => "11101010",
                     11850 => "01000001",
                     11851 => "00100111",
                     11852 => "10110010",
                     11853 => "10110011",
                     11854 => "01000010",
                     11855 => "00010110",
                     11856 => "11010100",
                     11857 => "01001010",
                     11858 => "01000010",
                     11859 => "10100101",
                     11860 => "01010001",
                     11861 => "10100111",
                     11862 => "00110001",
                     11863 => "00100111",
                     11864 => "11010011",
                     11865 => "00001000",
                     11866 => "11100010",
                     11867 => "00010110",
                     11868 => "01100100",
                     11869 => "00101100",
                     11870 => "00000100",
                     11871 => "00111000",
                     11872 => "01000010",
                     11873 => "01110110",
                     11874 => "01100100",
                     11875 => "10001000",
                     11876 => "01100010",
                     11877 => "11011110",
                     11878 => "00000111",
                     11879 => "11111110",
                     11880 => "00000001",
                     11881 => "00001101",
                     11882 => "11001001",
                     11883 => "00100011",
                     11884 => "00110010",
                     11885 => "00110001",
                     11886 => "01010001",
                     11887 => "10011000",
                     11888 => "01010010",
                     11889 => "00001101",
                     11890 => "11001001",
                     11891 => "01011001",
                     11892 => "01000010",
                     11893 => "01100011",
                     11894 => "01010011",
                     11895 => "01100111",
                     11896 => "00110001",
                     11897 => "00010100",
                     11898 => "11000010",
                     11899 => "00110110",
                     11900 => "00110001",
                     11901 => "10000111",
                     11902 => "01010011",
                     11903 => "00010111",
                     11904 => "11100011",
                     11905 => "00101001",
                     11906 => "01100001",
                     11907 => "00110000",
                     11908 => "01100010",
                     11909 => "00111100",
                     11910 => "00001000",
                     11911 => "01000010",
                     11912 => "00110111",
                     11913 => "01011001",
                     11914 => "01000000",
                     11915 => "01101010",
                     11916 => "01000010",
                     11917 => "10011001",
                     11918 => "01000000",
                     11919 => "11001001",
                     11920 => "01100001",
                     11921 => "11010111",
                     11922 => "01100011",
                     11923 => "00111001",
                     11924 => "11010001",
                     11925 => "01011000",
                     11926 => "01010010",
                     11927 => "11000011",
                     11928 => "01100111",
                     11929 => "11010011",
                     11930 => "00110001",
                     11931 => "11011100",
                     11932 => "00000110",
                     11933 => "11110111",
                     11934 => "01000010",
                     11935 => "11111010",
                     11936 => "01000010",
                     11937 => "00100011",
                     11938 => "10110001",
                     11939 => "01000011",
                     11940 => "01100111",
                     11941 => "11000011",
                     11942 => "00110100",
                     11943 => "11000111",
                     11944 => "00110100",
                     11945 => "11010001",
                     11946 => "01010001",
                     11947 => "01000011",
                     11948 => "10110011",
                     11949 => "01000111",
                     11950 => "00110011",
                     11951 => "10011010",
                     11952 => "00110000",
                     11953 => "10101001",
                     11954 => "01100001",
                     11955 => "10111000",
                     11956 => "01100010",
                     11957 => "10111110",
                     11958 => "00001011",
                     11959 => "11001110",
                     11960 => "00001111",
                     11961 => "11010101",
                     11962 => "00001001",
                     11963 => "00001101",
                     11964 => "11001010",
                     11965 => "01111101",
                     11966 => "01000111",
                     11967 => "11111101",
                     11968 => "01001001",
                     11969 => "00001111",
                     11970 => "00011110",
                     11971 => "00000001",
                     11972 => "00111001",
                     11973 => "01110011",
                     11974 => "01011110",
                     11975 => "00000111",
                     11976 => "10101110",
                     11977 => "00001011",
                     11978 => "00011110",
                     11979 => "10000010",
                     11980 => "01101110",
                     11981 => "10001000",
                     11982 => "10011110",
                     11983 => "00000010",
                     11984 => "00001101",
                     11985 => "00000100",
                     11986 => "00101110",
                     11987 => "00001011",
                     11988 => "00111110",
                     11989 => "00001111",
                     11990 => "01000101",
                     11991 => "00001001",
                     11992 => "11101101",
                     11993 => "01000111",
                     11994 => "11111101",
                     11995 => "11111111",
                     11996 => "10101101",
                     11997 => "01110010",
                     11998 => "00000111",
                     11999 => "00100000",
                     12000 => "00000100",
                     12001 => "10001110",
                     12002 => "11100100",
                     12003 => "10001111",
                     12004 => "01100111",
                     12005 => "10000101",
                     12006 => "01110001",
                     12007 => "10010000",
                     12008 => "11101010",
                     12009 => "10101110",
                     12010 => "10101110",
                     12011 => "01010011",
                     12012 => "00000111",
                     12013 => "10111101",
                     12014 => "11111100",
                     12015 => "00000110",
                     12016 => "10001101",
                     12017 => "11111100",
                     12018 => "00000110",
                     12019 => "00100000",
                     12020 => "01001010",
                     12021 => "10110000",
                     12022 => "10101101",
                     12023 => "01110010",
                     12024 => "00000111",
                     12025 => "11001001",
                     12026 => "00000011",
                     12027 => "10110000",
                     12028 => "00000001",
                     12029 => "01100000",
                     12030 => "00100000",
                     12031 => "00100100",
                     12032 => "10110110",
                     12033 => "10100010",
                     12034 => "00000000",
                     12035 => "10000110",
                     12036 => "00001000",
                     12037 => "00100000",
                     12038 => "01001101",
                     12039 => "11000000",
                     12040 => "00100000",
                     12041 => "11000011",
                     12042 => "10000100",
                     12043 => "11101000",
                     12044 => "11100000",
                     12045 => "00000110",
                     12046 => "11010000",
                     12047 => "11110011",
                     12048 => "00100000",
                     12049 => "10000111",
                     12050 => "11110001",
                     12051 => "00100000",
                     12052 => "00110001",
                     12053 => "11110001",
                     12054 => "00100000",
                     12055 => "11110000",
                     12056 => "11101110",
                     12057 => "00100000",
                     12058 => "11011001",
                     12059 => "10111110",
                     12060 => "10100010",
                     12061 => "00000001",
                     12062 => "10000110",
                     12063 => "00001000",
                     12064 => "00100000",
                     12065 => "01110101",
                     12066 => "10111110",
                     12067 => "11001010",
                     12068 => "10000110",
                     12069 => "00001000",
                     12070 => "00100000",
                     12071 => "01110101",
                     12072 => "10111110",
                     12073 => "00100000",
                     12074 => "10011011",
                     12075 => "10111011",
                     12076 => "00100000",
                     12077 => "11000001",
                     12078 => "10111001",
                     12079 => "00100000",
                     12080 => "10111000",
                     12081 => "10110111",
                     12082 => "00100000",
                     12083 => "01010101",
                     12084 => "10111000",
                     12085 => "00100000",
                     12086 => "01001111",
                     12087 => "10110111",
                     12088 => "00100000",
                     12089 => "11100001",
                     12090 => "10001001",
                     12091 => "10100101",
                     12092 => "10110101",
                     12093 => "11001001",
                     12094 => "00000010",
                     12095 => "00010000",
                     12096 => "00010001",
                     12097 => "10101101",
                     12098 => "10011111",
                     12099 => "00000111",
                     12100 => "11110000",
                     12101 => "00011110",
                     12102 => "11001001",
                     12103 => "00000100",
                     12104 => "11010000",
                     12105 => "00001000",
                     12106 => "10101101",
                     12107 => "01111111",
                     12108 => "00000111",
                     12109 => "11010000",
                     12110 => "00000011",
                     12111 => "00100000",
                     12112 => "11101101",
                     12113 => "10010000",
                     12114 => "10101100",
                     12115 => "10011111",
                     12116 => "00000111",
                     12117 => "10100101",
                     12118 => "00001001",
                     12119 => "11000000",
                     12120 => "00001000",
                     12121 => "10110000",
                     12122 => "00000010",
                     12123 => "01001010",
                     12124 => "01001010",
                     12125 => "01001010",
                     12126 => "00100000",
                     12127 => "10001000",
                     12128 => "10110010",
                     12129 => "01001100",
                     12130 => "01100111",
                     12131 => "10101111",
                     12132 => "00100000",
                     12133 => "10011010",
                     12134 => "10110010",
                     12135 => "10100101",
                     12136 => "00001010",
                     12137 => "10000101",
                     12138 => "00001101",
                     12139 => "10101001",
                     12140 => "00000000",
                     12141 => "10000101",
                     12142 => "00001100",
                     12143 => "10101101",
                     12144 => "01110011",
                     12145 => "00000111",
                     12146 => "11001001",
                     12147 => "00000110",
                     12148 => "11110000",
                     12149 => "00011100",
                     12150 => "10101101",
                     12151 => "00011111",
                     12152 => "00000111",
                     12153 => "11010000",
                     12154 => "00010100",
                     12155 => "10101101",
                     12156 => "00111101",
                     12157 => "00000111",
                     12158 => "11001001",
                     12159 => "00100000",
                     12160 => "00110000",
                     12161 => "00010000",
                     12162 => "10101101",
                     12163 => "00111101",
                     12164 => "00000111",
                     12165 => "11101001",
                     12166 => "00100000",
                     12167 => "10001101",
                     12168 => "00111101",
                     12169 => "00000111",
                     12170 => "10101001",
                     12171 => "00000000",
                     12172 => "10001101",
                     12173 => "01000000",
                     12174 => "00000011",
                     12175 => "00100000",
                     12176 => "10110000",
                     12177 => "10010010",
                     12178 => "01100000",
                     12179 => "10101101",
                     12180 => "11111111",
                     12181 => "00000110",
                     12182 => "00011000",
                     12183 => "01101101",
                     12184 => "10100001",
                     12185 => "00000011",
                     12186 => "10001101",
                     12187 => "11111111",
                     12188 => "00000110",
                     12189 => "10101101",
                     12190 => "00100011",
                     12191 => "00000111",
                     12192 => "11010000",
                     12193 => "01011001",
                     12194 => "10101101",
                     12195 => "01010101",
                     12196 => "00000111",
                     12197 => "11001001",
                     12198 => "01010000",
                     12199 => "10010000",
                     12200 => "01010010",
                     12201 => "10101101",
                     12202 => "10000101",
                     12203 => "00000111",
                     12204 => "11010000",
                     12205 => "01001101",
                     12206 => "10101100",
                     12207 => "11111111",
                     12208 => "00000110",
                     12209 => "10001000",
                     12210 => "00110000",
                     12211 => "01000111",
                     12212 => "11001000",
                     12213 => "11000000",
                     12214 => "00000010",
                     12215 => "10010000",
                     12216 => "00000001",
                     12217 => "10001000",
                     12218 => "10101101",
                     12219 => "01010101",
                     12220 => "00000111",
                     12221 => "11001001",
                     12222 => "01110000",
                     12223 => "10010000",
                     12224 => "00000011",
                     12225 => "10101100",
                     12226 => "11111111",
                     12227 => "00000110",
                     12228 => "10011000",
                     12229 => "10001101",
                     12230 => "01110101",
                     12231 => "00000111",
                     12232 => "00011000",
                     12233 => "01101101",
                     12234 => "00111101",
                     12235 => "00000111",
                     12236 => "10001101",
                     12237 => "00111101",
                     12238 => "00000111",
                     12239 => "10011000",
                     12240 => "00011000",
                     12241 => "01101101",
                     12242 => "00011100",
                     12243 => "00000111",
                     12244 => "10001101",
                     12245 => "00011100",
                     12246 => "00000111",
                     12247 => "10001101",
                     12248 => "00111111",
                     12249 => "00000111",
                     12250 => "10101101",
                     12251 => "00011010",
                     12252 => "00000111",
                     12253 => "01101001",
                     12254 => "00000000",
                     12255 => "10001101",
                     12256 => "00011010",
                     12257 => "00000111",
                     12258 => "00101001",
                     12259 => "00000001",
                     12260 => "10000101",
                     12261 => "00000000",
                     12262 => "10101101",
                     12263 => "01111000",
                     12264 => "00000111",
                     12265 => "00101001",
                     12266 => "11111110",
                     12267 => "00000101",
                     12268 => "00000000",
                     12269 => "10001101",
                     12270 => "01111000",
                     12271 => "00000111",
                     12272 => "00100000",
                     12273 => "00111000",
                     12274 => "10110000",
                     12275 => "10101001",
                     12276 => "00001000",
                     12277 => "10001101",
                     12278 => "10010101",
                     12279 => "00000111",
                     12280 => "01001100",
                     12281 => "00000000",
                     12282 => "10110000",
                     12283 => "10101001",
                     12284 => "00000000",
                     12285 => "10001101",
                     12286 => "01110101",
                     12287 => "00000111",
                     12288 => "10100010",
                     12289 => "00000000",
                     12290 => "00100000",
                     12291 => "11111101",
                     12292 => "11110001",
                     12293 => "10000101",
                     12294 => "00000000",
                     12295 => "10100000",
                     12296 => "00000000",
                     12297 => "00001010",
                     12298 => "10110000",
                     12299 => "00000111",
                     12300 => "11001000",
                     12301 => "10100101",
                     12302 => "00000000",
                     12303 => "00101001",
                     12304 => "00100000",
                     12305 => "11110000",
                     12306 => "00011011",
                     12307 => "10111001",
                     12308 => "00011100",
                     12309 => "00000111",
                     12310 => "00111000",
                     12311 => "11111001",
                     12312 => "00110100",
                     12313 => "10110000",
                     12314 => "10000101",
                     12315 => "10000110",
                     12316 => "10111001",
                     12317 => "00011010",
                     12318 => "00000111",
                     12319 => "11101001",
                     12320 => "00000000",
                     12321 => "10000101",
                     12322 => "01101101",
                     12323 => "10100101",
                     12324 => "00001100",
                     12325 => "11011001",
                     12326 => "00110110",
                     12327 => "10110000",
                     12328 => "11110000",
                     12329 => "00000100",
                     12330 => "10101001",
                     12331 => "00000000",
                     12332 => "10000101",
                     12333 => "01010111",
                     12334 => "10101001",
                     12335 => "00000000",
                     12336 => "10001101",
                     12337 => "10100001",
                     12338 => "00000011",
                     12339 => "01100000",
                     12340 => "00000000",
                     12341 => "00010000",
                     12342 => "00000001",
                     12343 => "00000010",
                     12344 => "10101101",
                     12345 => "00011100",
                     12346 => "00000111",
                     12347 => "00011000",
                     12348 => "01101001",
                     12349 => "11111111",
                     12350 => "10001101",
                     12351 => "00011101",
                     12352 => "00000111",
                     12353 => "10101101",
                     12354 => "00011010",
                     12355 => "00000111",
                     12356 => "01101001",
                     12357 => "00000000",
                     12358 => "10001101",
                     12359 => "00011011",
                     12360 => "00000111",
                     12361 => "01100000",
                     12362 => "10100101",
                     12363 => "00001110",
                     12364 => "00100000",
                     12365 => "00000100",
                     12366 => "10001110",
                     12367 => "00110001",
                     12368 => "10010001",
                     12369 => "11000111",
                     12370 => "10110001",
                     12371 => "00000110",
                     12372 => "10110010",
                     12373 => "11100101",
                     12374 => "10110001",
                     12375 => "10100100",
                     12376 => "10110010",
                     12377 => "11001010",
                     12378 => "10110010",
                     12379 => "11001101",
                     12380 => "10010001",
                     12381 => "01101001",
                     12382 => "10110000",
                     12383 => "11101001",
                     12384 => "10110000",
                     12385 => "00110011",
                     12386 => "10110010",
                     12387 => "01000101",
                     12388 => "10110010",
                     12389 => "01101001",
                     12390 => "10110010",
                     12391 => "01111101",
                     12392 => "10110010",
                     12393 => "10101101",
                     12394 => "01010010",
                     12395 => "00000111",
                     12396 => "11001001",
                     12397 => "00000010",
                     12398 => "11110000",
                     12399 => "00101011",
                     12400 => "10101001",
                     12401 => "00000000",
                     12402 => "10100100",
                     12403 => "11001110",
                     12404 => "11000000",
                     12405 => "00110000",
                     12406 => "10010000",
                     12407 => "01101110",
                     12408 => "10101101",
                     12409 => "00010000",
                     12410 => "00000111",
                     12411 => "11001001",
                     12412 => "00000110",
                     12413 => "11110000",
                     12414 => "00000100",
                     12415 => "11001001",
                     12416 => "00000111",
                     12417 => "11010000",
                     12418 => "01010000",
                     12419 => "10101101",
                     12420 => "11000100",
                     12421 => "00000011",
                     12422 => "11010000",
                     12423 => "00000101",
                     12424 => "10101001",
                     12425 => "00000001",
                     12426 => "01001100",
                     12427 => "11100110",
                     12428 => "10110000",
                     12429 => "00100000",
                     12430 => "00011111",
                     12431 => "10110010",
                     12432 => "11001110",
                     12433 => "11011110",
                     12434 => "00000110",
                     12435 => "11010000",
                     12436 => "01010000",
                     12437 => "11101110",
                     12438 => "01101001",
                     12439 => "00000111",
                     12440 => "01001100",
                     12441 => "00010101",
                     12442 => "10110011",
                     12443 => "10101101",
                     12444 => "01011000",
                     12445 => "00000111",
                     12446 => "11010000",
                     12447 => "00001100",
                     12448 => "10101001",
                     12449 => "11111111",
                     12450 => "00100000",
                     12451 => "00000000",
                     12452 => "10110010",
                     12453 => "10100101",
                     12454 => "11001110",
                     12455 => "11001001",
                     12456 => "10010001",
                     12457 => "10010000",
                     12458 => "00101000",
                     12459 => "01100000",
                     12460 => "10101101",
                     12461 => "10011001",
                     12462 => "00000011",
                     12463 => "11001001",
                     12464 => "01100000",
                     12465 => "11010000",
                     12466 => "00110010",
                     12467 => "10100101",
                     12468 => "11001110",
                     12469 => "11001001",
                     12470 => "10011001",
                     12471 => "10100000",
                     12472 => "00000000",
                     12473 => "10101001",
                     12474 => "00000001",
                     12475 => "10010000",
                     12476 => "00001010",
                     12477 => "10101001",
                     12478 => "00000011",
                     12479 => "10000101",
                     12480 => "00011101",
                     12481 => "11001000",
                     12482 => "10101001",
                     12483 => "00001000",
                     12484 => "10001101",
                     12485 => "10110100",
                     12486 => "00000101",
                     12487 => "10001100",
                     12488 => "00010110",
                     12489 => "00000111",
                     12490 => "00100000",
                     12491 => "11100110",
                     12492 => "10110000",
                     12493 => "10100101",
                     12494 => "10000110",
                     12495 => "11001001",
                     12496 => "01001000",
                     12497 => "10010000",
                     12498 => "00010010",
                     12499 => "10101001",
                     12500 => "00001000",
                     12501 => "10000101",
                     12502 => "00001110",
                     12503 => "10101001",
                     12504 => "00000001",
                     12505 => "10000101",
                     12506 => "00110011",
                     12507 => "01001010",
                     12508 => "10001101",
                     12509 => "01010010",
                     12510 => "00000111",
                     12511 => "10001101",
                     12512 => "00010110",
                     12513 => "00000111",
                     12514 => "10001101",
                     12515 => "01011000",
                     12516 => "00000111",
                     12517 => "01100000",
                     12518 => "10001101",
                     12519 => "11111100",
                     12520 => "00000110",
                     12521 => "10100101",
                     12522 => "00001110",
                     12523 => "11001001",
                     12524 => "00001011",
                     12525 => "11110000",
                     12526 => "00111100",
                     12527 => "10101101",
                     12528 => "01001110",
                     12529 => "00000111",
                     12530 => "11010000",
                     12531 => "00010000",
                     12532 => "10100100",
                     12533 => "10110101",
                     12534 => "10001000",
                     12535 => "11010000",
                     12536 => "00000110",
                     12537 => "10100101",
                     12538 => "11001110",
                     12539 => "11001001",
                     12540 => "11010000",
                     12541 => "10010000",
                     12542 => "00000101",
                     12543 => "10101001",
                     12544 => "00000000",
                     12545 => "10001101",
                     12546 => "11111100",
                     12547 => "00000110",
                     12548 => "10101101",
                     12549 => "11111100",
                     12550 => "00000110",
                     12551 => "00101001",
                     12552 => "11000000",
                     12553 => "10000101",
                     12554 => "00001010",
                     12555 => "10101101",
                     12556 => "11111100",
                     12557 => "00000110",
                     12558 => "00101001",
                     12559 => "00000011",
                     12560 => "10000101",
                     12561 => "00001100",
                     12562 => "10101101",
                     12563 => "11111100",
                     12564 => "00000110",
                     12565 => "00101001",
                     12566 => "00001100",
                     12567 => "10000101",
                     12568 => "00001011",
                     12569 => "00101001",
                     12570 => "00000100",
                     12571 => "11110000",
                     12572 => "00001110",
                     12573 => "10100101",
                     12574 => "00011101",
                     12575 => "11010000",
                     12576 => "00001010",
                     12577 => "10100100",
                     12578 => "00001100",
                     12579 => "11110000",
                     12580 => "00000110",
                     12581 => "10101001",
                     12582 => "00000000",
                     12583 => "10000101",
                     12584 => "00001100",
                     12585 => "10000101",
                     12586 => "00001011",
                     12587 => "00100000",
                     12588 => "00101001",
                     12589 => "10110011",
                     12590 => "10100000",
                     12591 => "00000001",
                     12592 => "10101101",
                     12593 => "01010100",
                     12594 => "00000111",
                     12595 => "11010000",
                     12596 => "00001001",
                     12597 => "10100000",
                     12598 => "00000000",
                     12599 => "10101101",
                     12600 => "00010100",
                     12601 => "00000111",
                     12602 => "11110000",
                     12603 => "00000010",
                     12604 => "10100000",
                     12605 => "00000010",
                     12606 => "10001100",
                     12607 => "10011001",
                     12608 => "00000100",
                     12609 => "10101001",
                     12610 => "00000001",
                     12611 => "10100100",
                     12612 => "01010111",
                     12613 => "11110000",
                     12614 => "00000101",
                     12615 => "00010000",
                     12616 => "00000001",
                     12617 => "00001010",
                     12618 => "10000101",
                     12619 => "01000101",
                     12620 => "00100000",
                     12621 => "10010011",
                     12622 => "10101111",
                     12623 => "00100000",
                     12624 => "10000111",
                     12625 => "11110001",
                     12626 => "00100000",
                     12627 => "00110001",
                     12628 => "11110001",
                     12629 => "10100010",
                     12630 => "00000000",
                     12631 => "00100000",
                     12632 => "10100100",
                     12633 => "11100010",
                     12634 => "00100000",
                     12635 => "01100110",
                     12636 => "11011100",
                     12637 => "10100101",
                     12638 => "11001110",
                     12639 => "11001001",
                     12640 => "01000000",
                     12641 => "10010000",
                     12642 => "00010110",
                     12643 => "10100101",
                     12644 => "00001110",
                     12645 => "11001001",
                     12646 => "00000101",
                     12647 => "11110000",
                     12648 => "00010000",
                     12649 => "11001001",
                     12650 => "00000111",
                     12651 => "11110000",
                     12652 => "00001100",
                     12653 => "11001001",
                     12654 => "00000100",
                     12655 => "10010000",
                     12656 => "00001000",
                     12657 => "10101101",
                     12658 => "11000100",
                     12659 => "00000011",
                     12660 => "00101001",
                     12661 => "11011111",
                     12662 => "10001101",
                     12663 => "11000100",
                     12664 => "00000011",
                     12665 => "10100101",
                     12666 => "10110101",
                     12667 => "11001001",
                     12668 => "00000010",
                     12669 => "00110000",
                     12670 => "00111011",
                     12671 => "10100010",
                     12672 => "00000001",
                     12673 => "10001110",
                     12674 => "00100011",
                     12675 => "00000111",
                     12676 => "10100000",
                     12677 => "00000100",
                     12678 => "10000100",
                     12679 => "00000111",
                     12680 => "10100010",
                     12681 => "00000000",
                     12682 => "10101100",
                     12683 => "01011001",
                     12684 => "00000111",
                     12685 => "11010000",
                     12686 => "00000101",
                     12687 => "10101100",
                     12688 => "01000011",
                     12689 => "00000111",
                     12690 => "11010000",
                     12691 => "00010110",
                     12692 => "11101000",
                     12693 => "10100100",
                     12694 => "00001110",
                     12695 => "11000000",
                     12696 => "00001011",
                     12697 => "11110000",
                     12698 => "00001111",
                     12699 => "10101100",
                     12700 => "00010010",
                     12701 => "00000111",
                     12702 => "11010000",
                     12703 => "00000110",
                     12704 => "11001000",
                     12705 => "10000100",
                     12706 => "11111100",
                     12707 => "10001100",
                     12708 => "00010010",
                     12709 => "00000111",
                     12710 => "10100000",
                     12711 => "00000110",
                     12712 => "10000100",
                     12713 => "00000111",
                     12714 => "11000101",
                     12715 => "00000111",
                     12716 => "00110000",
                     12717 => "00001100",
                     12718 => "11001010",
                     12719 => "00110000",
                     12720 => "00001010",
                     12721 => "10101100",
                     12722 => "10110001",
                     12723 => "00000111",
                     12724 => "11010000",
                     12725 => "00000100",
                     12726 => "10101001",
                     12727 => "00000110",
                     12728 => "10000101",
                     12729 => "00001110",
                     12730 => "01100000",
                     12731 => "10101001",
                     12732 => "00000000",
                     12733 => "10001101",
                     12734 => "01011000",
                     12735 => "00000111",
                     12736 => "00100000",
                     12737 => "11011101",
                     12738 => "10110001",
                     12739 => "11101110",
                     12740 => "01010010",
                     12741 => "00000111",
                     12742 => "01100000",
                     12743 => "10100101",
                     12744 => "10110101",
                     12745 => "11010000",
                     12746 => "00000110",
                     12747 => "10100101",
                     12748 => "11001110",
                     12749 => "11001001",
                     12750 => "11100100",
                     12751 => "10010000",
                     12752 => "00001100",
                     12753 => "10101001",
                     12754 => "00001000",
                     12755 => "10001101",
                     12756 => "01011000",
                     12757 => "00000111",
                     12758 => "10100000",
                     12759 => "00000011",
                     12760 => "10000100",
                     12761 => "00011101",
                     12762 => "01001100",
                     12763 => "11100110",
                     12764 => "10110000",
                     12765 => "10101001",
                     12766 => "00000010",
                     12767 => "10001101",
                     12768 => "01010010",
                     12769 => "00000111",
                     12770 => "01001100",
                     12771 => "00010011",
                     12772 => "10110010",
                     12773 => "10101001",
                     12774 => "00000001",
                     12775 => "00100000",
                     12776 => "00000000",
                     12777 => "10110010",
                     12778 => "00100000",
                     12779 => "10010011",
                     12780 => "10101111",
                     12781 => "10100000",
                     12782 => "00000000",
                     12783 => "10101101",
                     12784 => "11010110",
                     12785 => "00000110",
                     12786 => "11010000",
                     12787 => "00010111",
                     12788 => "11001000",
                     12789 => "10101101",
                     12790 => "01001110",
                     12791 => "00000111",
                     12792 => "11001001",
                     12793 => "00000011",
                     12794 => "11010000",
                     12795 => "00001111",
                     12796 => "11001000",
                     12797 => "01001100",
                     12798 => "00001011",
                     12799 => "10110010",
                     12800 => "00011000",
                     12801 => "01100101",
                     12802 => "11001110",
                     12803 => "10000101",
                     12804 => "11001110",
                     12805 => "01100000",
                     12806 => "00100000",
                     12807 => "00011111",
                     12808 => "10110010",
                     12809 => "10100000",
                     12810 => "00000010",
                     12811 => "11001110",
                     12812 => "11011110",
                     12813 => "00000110",
                     12814 => "11010000",
                     12815 => "00001110",
                     12816 => "10001100",
                     12817 => "01010010",
                     12818 => "00000111",
                     12819 => "11101110",
                     12820 => "01110100",
                     12821 => "00000111",
                     12822 => "10101001",
                     12823 => "00000000",
                     12824 => "10001101",
                     12825 => "01110010",
                     12826 => "00000111",
                     12827 => "10001101",
                     12828 => "00100010",
                     12829 => "00000111",
                     12830 => "01100000",
                     12831 => "10101001",
                     12832 => "00001000",
                     12833 => "10000101",
                     12834 => "01010111",
                     12835 => "10100000",
                     12836 => "00000001",
                     12837 => "10100101",
                     12838 => "10000110",
                     12839 => "00101001",
                     12840 => "00001111",
                     12841 => "11010000",
                     12842 => "00000011",
                     12843 => "10000101",
                     12844 => "01010111",
                     12845 => "10101000",
                     12846 => "10011000",
                     12847 => "00100000",
                     12848 => "11100110",
                     12849 => "10110000",
                     12850 => "01100000",
                     12851 => "10101101",
                     12852 => "01000111",
                     12853 => "00000111",
                     12854 => "11001001",
                     12855 => "11111000",
                     12856 => "11010000",
                     12857 => "00000011",
                     12858 => "01001100",
                     12859 => "01010101",
                     12860 => "10110010",
                     12861 => "11001001",
                     12862 => "11000100",
                     12863 => "11010000",
                     12864 => "00000011",
                     12865 => "00100000",
                     12866 => "01110011",
                     12867 => "10110010",
                     12868 => "01100000",
                     12869 => "10101101",
                     12870 => "01000111",
                     12871 => "00000111",
                     12872 => "11001001",
                     12873 => "11110000",
                     12874 => "10110000",
                     12875 => "00000111",
                     12876 => "11001001",
                     12877 => "11001000",
                     12878 => "11110000",
                     12879 => "00100011",
                     12880 => "01001100",
                     12881 => "11101001",
                     12882 => "10110000",
                     12883 => "11010000",
                     12884 => "00010011",
                     12885 => "10101100",
                     12886 => "00001011",
                     12887 => "00000111",
                     12888 => "11010000",
                     12889 => "00001110",
                     12890 => "10001100",
                     12891 => "00001101",
                     12892 => "00000111",
                     12893 => "11101110",
                     12894 => "00001011",
                     12895 => "00000111",
                     12896 => "10101101",
                     12897 => "01010100",
                     12898 => "00000111",
                     12899 => "01001001",
                     12900 => "00000001",
                     12901 => "10001101",
                     12902 => "01010100",
                     12903 => "00000111",
                     12904 => "01100000",
                     12905 => "10101101",
                     12906 => "01000111",
                     12907 => "00000111",
                     12908 => "11001001",
                     12909 => "11110000",
                     12910 => "10110000",
                     12911 => "00110011",
                     12912 => "01001100",
                     12913 => "11101001",
                     12914 => "10110000",
                     12915 => "10101001",
                     12916 => "00000000",
                     12917 => "10001101",
                     12918 => "01000111",
                     12919 => "00000111",
                     12920 => "10101001",
                     12921 => "00001000",
                     12922 => "10000101",
                     12923 => "00001110",
                     12924 => "01100000",
                     12925 => "10101101",
                     12926 => "01000111",
                     12927 => "00000111",
                     12928 => "11001001",
                     12929 => "11000000",
                     12930 => "11110000",
                     12931 => "00010011",
                     12932 => "10100101",
                     12933 => "00001001",
                     12934 => "01001010",
                     12935 => "01001010",
                     12936 => "00101001",
                     12937 => "00000011",
                     12938 => "10000101",
                     12939 => "00000000",
                     12940 => "10101101",
                     12941 => "11000100",
                     12942 => "00000011",
                     12943 => "00101001",
                     12944 => "11111100",
                     12945 => "00000101",
                     12946 => "00000000",
                     12947 => "10001101",
                     12948 => "11000100",
                     12949 => "00000011",
                     12950 => "01100000",
                     12951 => "00100000",
                     12952 => "01110011",
                     12953 => "10110010",
                     12954 => "10101101",
                     12955 => "11000100",
                     12956 => "00000011",
                     12957 => "00101001",
                     12958 => "11111100",
                     12959 => "10001101",
                     12960 => "11000100",
                     12961 => "00000011",
                     12962 => "01100000",
                     12963 => "01100000",
                     12964 => "10100101",
                     12965 => "00011011",
                     12966 => "11001001",
                     12967 => "00110000",
                     12968 => "11010000",
                     12969 => "00010101",
                     12970 => "10101101",
                     12971 => "00010011",
                     12972 => "00000111",
                     12973 => "10000101",
                     12974 => "11111111",
                     12975 => "10101001",
                     12976 => "00000000",
                     12977 => "10001101",
                     12978 => "00010011",
                     12979 => "00000111",
                     12980 => "10100100",
                     12981 => "11001110",
                     12982 => "11000000",
                     12983 => "10011110",
                     12984 => "10110000",
                     12985 => "00000010",
                     12986 => "10101001",
                     12987 => "00000100",
                     12988 => "01001100",
                     12989 => "11100110",
                     12990 => "10110000",
                     12991 => "11100110",
                     12992 => "00001110",
                     12993 => "01100000",
                     12994 => "00010101",
                     12995 => "00100011",
                     12996 => "00010110",
                     12997 => "00011011",
                     12998 => "00010111",
                     12999 => "00011000",
                     13000 => "00100011",
                     13001 => "01100011",
                     13002 => "10101001",
                     13003 => "00000001",
                     13004 => "00100000",
                     13005 => "11100110",
                     13006 => "10110000",
                     13007 => "10100101",
                     13008 => "11001110",
                     13009 => "11001001",
                     13010 => "10101110",
                     13011 => "10010000",
                     13012 => "00001110",
                     13013 => "10101101",
                     13014 => "00100011",
                     13015 => "00000111",
                     13016 => "11110000",
                     13017 => "00001001",
                     13018 => "10101001",
                     13019 => "00100000",
                     13020 => "10000101",
                     13021 => "11111100",
                     13022 => "10101001",
                     13023 => "00000000",
                     13024 => "10001101",
                     13025 => "00100011",
                     13026 => "00000111",
                     13027 => "10101101",
                     13028 => "10010000",
                     13029 => "00000100",
                     13030 => "01001010",
                     13031 => "10110000",
                     13032 => "00001101",
                     13033 => "10101101",
                     13034 => "01000110",
                     13035 => "00000111",
                     13036 => "11010000",
                     13037 => "00000011",
                     13038 => "11101110",
                     13039 => "01000110",
                     13040 => "00000111",
                     13041 => "10101001",
                     13042 => "00100000",
                     13043 => "10001101",
                     13044 => "11000100",
                     13045 => "00000011",
                     13046 => "10101101",
                     13047 => "01000110",
                     13048 => "00000111",
                     13049 => "11001001",
                     13050 => "00000101",
                     13051 => "11010000",
                     13052 => "00101011",
                     13053 => "11101110",
                     13054 => "01011100",
                     13055 => "00000111",
                     13056 => "10101101",
                     13057 => "01011100",
                     13058 => "00000111",
                     13059 => "11001001",
                     13060 => "00000011",
                     13061 => "11010000",
                     13062 => "00001110",
                     13063 => "10101100",
                     13064 => "01011111",
                     13065 => "00000111",
                     13066 => "10101101",
                     13067 => "01001000",
                     13068 => "00000111",
                     13069 => "11011001",
                     13070 => "11000010",
                     13071 => "10110010",
                     13072 => "10010000",
                     13073 => "00000011",
                     13074 => "11101110",
                     13075 => "01011101",
                     13076 => "00000111",
                     13077 => "11101110",
                     13078 => "01100000",
                     13079 => "00000111",
                     13080 => "00100000",
                     13081 => "00000011",
                     13082 => "10011100",
                     13083 => "11101110",
                     13084 => "01010111",
                     13085 => "00000111",
                     13086 => "00100000",
                     13087 => "00010011",
                     13088 => "10110010",
                     13089 => "10001101",
                     13090 => "01011011",
                     13091 => "00000111",
                     13092 => "10101001",
                     13093 => "10000000",
                     13094 => "10000101",
                     13095 => "11111100",
                     13096 => "01100000",
                     13097 => "10101001",
                     13098 => "00000000",
                     13099 => "10101100",
                     13100 => "01010100",
                     13101 => "00000111",
                     13102 => "11010000",
                     13103 => "00001000",
                     13104 => "10100101",
                     13105 => "00011101",
                     13106 => "11010000",
                     13107 => "00000111",
                     13108 => "10100101",
                     13109 => "00001011",
                     13110 => "00101001",
                     13111 => "00000100",
                     13112 => "10001101",
                     13113 => "00010100",
                     13114 => "00000111",
                     13115 => "00100000",
                     13116 => "01010000",
                     13117 => "10110100",
                     13118 => "10101101",
                     13119 => "00001011",
                     13120 => "00000111",
                     13121 => "11010000",
                     13122 => "00010110",
                     13123 => "10100101",
                     13124 => "00011101",
                     13125 => "11001001",
                     13126 => "00000011",
                     13127 => "11110000",
                     13128 => "00000101",
                     13129 => "10100000",
                     13130 => "00011000",
                     13131 => "10001100",
                     13132 => "10001001",
                     13133 => "00000111",
                     13134 => "00100000",
                     13135 => "00000100",
                     13136 => "10001110",
                     13137 => "01011010",
                     13138 => "10110011",
                     13139 => "01110110",
                     13140 => "10110011",
                     13141 => "01101101",
                     13142 => "10110011",
                     13143 => "11001111",
                     13144 => "10110011",
                     13145 => "01100000",
                     13146 => "00100000",
                     13147 => "10001111",
                     13148 => "10110101",
                     13149 => "10100101",
                     13150 => "00001100",
                     13151 => "11110000",
                     13152 => "00000010",
                     13153 => "10000101",
                     13154 => "00110011",
                     13155 => "00100000",
                     13156 => "11001100",
                     13157 => "10110101",
                     13158 => "00100000",
                     13159 => "00001110",
                     13160 => "10111111",
                     13161 => "10001101",
                     13162 => "11111111",
                     13163 => "00000110",
                     13164 => "01100000",
                     13165 => "10101101",
                     13166 => "00001010",
                     13167 => "00000111",
                     13168 => "10001101",
                     13169 => "00001001",
                     13170 => "00000111",
                     13171 => "01001100",
                     13172 => "10101100",
                     13173 => "10110011",
                     13174 => "10100100",
                     13175 => "10011111",
                     13176 => "00010000",
                     13177 => "00010011",
                     13178 => "10100101",
                     13179 => "00001010",
                     13180 => "00101001",
                     13181 => "10000000",
                     13182 => "00100101",
                     13183 => "00001101",
                     13184 => "11010000",
                     13185 => "00010001",
                     13186 => "10101101",
                     13187 => "00001000",
                     13188 => "00000111",
                     13189 => "00111000",
                     13190 => "11100101",
                     13191 => "11001110",
                     13192 => "11001101",
                     13193 => "00000110",
                     13194 => "00000111",
                     13195 => "10010000",
                     13196 => "00000110",
                     13197 => "10101101",
                     13198 => "00001010",
                     13199 => "00000111",
                     13200 => "10001101",
                     13201 => "00001001",
                     13202 => "00000111",
                     13203 => "10101101",
                     13204 => "00000100",
                     13205 => "00000111",
                     13206 => "11110000",
                     13207 => "00010100",
                     13208 => "00100000",
                     13209 => "10001111",
                     13210 => "10110101",
                     13211 => "10100101",
                     13212 => "11001110",
                     13213 => "11001001",
                     13214 => "00010100",
                     13215 => "10110000",
                     13216 => "00000101",
                     13217 => "10101001",
                     13218 => "00011000",
                     13219 => "10001101",
                     13220 => "00001001",
                     13221 => "00000111",
                     13222 => "10100101",
                     13223 => "00001100",
                     13224 => "11110000",
                     13225 => "00000010",
                     13226 => "10000101",
                     13227 => "00110011",
                     13228 => "10100101",
                     13229 => "00001100",
                     13230 => "11110000",
                     13231 => "00000011",
                     13232 => "00100000",
                     13233 => "11001100",
                     13234 => "10110101",
                     13235 => "00100000",
                     13236 => "00001110",
                     13237 => "10111111",
                     13238 => "10001101",
                     13239 => "11111111",
                     13240 => "00000110",
                     13241 => "10100101",
                     13242 => "00001110",
                     13243 => "11001001",
                     13244 => "00001011",
                     13245 => "11010000",
                     13246 => "00000101",
                     13247 => "10101001",
                     13248 => "00101000",
                     13249 => "10001101",
                     13250 => "00001001",
                     13251 => "00000111",
                     13252 => "01001100",
                     13253 => "01010010",
                     13254 => "10111111",
                     13255 => "00001110",
                     13256 => "00000100",
                     13257 => "11111100",
                     13258 => "11110010",
                     13259 => "00000000",
                     13260 => "00000000",
                     13261 => "11111111",
                     13262 => "11111111",
                     13263 => "10101101",
                     13264 => "00010110",
                     13265 => "00000100",
                     13266 => "00011000",
                     13267 => "01101101",
                     13268 => "00110011",
                     13269 => "00000100",
                     13270 => "10001101",
                     13271 => "00010110",
                     13272 => "00000100",
                     13273 => "10100000",
                     13274 => "00000000",
                     13275 => "10100101",
                     13276 => "10011111",
                     13277 => "00010000",
                     13278 => "00000001",
                     13279 => "10001000",
                     13280 => "10000100",
                     13281 => "00000000",
                     13282 => "01100101",
                     13283 => "11001110",
                     13284 => "10000101",
                     13285 => "11001110",
                     13286 => "10100101",
                     13287 => "10110101",
                     13288 => "01100101",
                     13289 => "00000000",
                     13290 => "10000101",
                     13291 => "10110101",
                     13292 => "10100101",
                     13293 => "00001100",
                     13294 => "00101101",
                     13295 => "10010000",
                     13296 => "00000100",
                     13297 => "11110000",
                     13298 => "00101101",
                     13299 => "10101100",
                     13300 => "10001001",
                     13301 => "00000111",
                     13302 => "11010000",
                     13303 => "00100111",
                     13304 => "10100000",
                     13305 => "00011000",
                     13306 => "10001100",
                     13307 => "10001001",
                     13308 => "00000111",
                     13309 => "10100010",
                     13310 => "00000000",
                     13311 => "10100100",
                     13312 => "00110011",
                     13313 => "01001010",
                     13314 => "10110000",
                     13315 => "00000010",
                     13316 => "11101000",
                     13317 => "11101000",
                     13318 => "10001000",
                     13319 => "11110000",
                     13320 => "00000001",
                     13321 => "11101000",
                     13322 => "10100101",
                     13323 => "10000110",
                     13324 => "00011000",
                     13325 => "01111101",
                     13326 => "11000111",
                     13327 => "10110011",
                     13328 => "10000101",
                     13329 => "10000110",
                     13330 => "10100101",
                     13331 => "01101101",
                     13332 => "01111101",
                     13333 => "11001011",
                     13334 => "10110011",
                     13335 => "10000101",
                     13336 => "01101101",
                     13337 => "10100101",
                     13338 => "00001100",
                     13339 => "01001001",
                     13340 => "00000011",
                     13341 => "10000101",
                     13342 => "00110011",
                     13343 => "01100000",
                     13344 => "10001101",
                     13345 => "10001001",
                     13346 => "00000111",
                     13347 => "01100000",
                     13348 => "00110000",
                     13349 => "00110000",
                     13350 => "00101101",
                     13351 => "00111000",
                     13352 => "00111000",
                     13353 => "00001101",
                     13354 => "00000100",
                     13355 => "10101000",
                     13356 => "10101000",
                     13357 => "10010000",
                     13358 => "11010000",
                     13359 => "11010000",
                     13360 => "00001010",
                     13361 => "00001001",
                     13362 => "11111011",
                     13363 => "11111011",
                     13364 => "11111011",
                     13365 => "11111010",
                     13366 => "11111010",
                     13367 => "11111110",
                     13368 => "11111111",
                     13369 => "00110100",
                     13370 => "00110100",
                     13371 => "00110100",
                     13372 => "00000000",
                     13373 => "00000000",
                     13374 => "10000000",
                     13375 => "00000000",
                     13376 => "11010000",
                     13377 => "11100100",
                     13378 => "11101101",
                     13379 => "00110000",
                     13380 => "00011100",
                     13381 => "00010011",
                     13382 => "00001110",
                     13383 => "11000000",
                     13384 => "00000000",
                     13385 => "10000000",
                     13386 => "00000000",
                     13387 => "11111111",
                     13388 => "00000001",
                     13389 => "00000000",
                     13390 => "00100000",
                     13391 => "11111111",
                     13392 => "10100101",
                     13393 => "00011101",
                     13394 => "11001001",
                     13395 => "00000011",
                     13396 => "11010000",
                     13397 => "00100011",
                     13398 => "10100000",
                     13399 => "00000000",
                     13400 => "10100101",
                     13401 => "00001011",
                     13402 => "00101101",
                     13403 => "10010000",
                     13404 => "00000100",
                     13405 => "11110000",
                     13406 => "00000110",
                     13407 => "11001000",
                     13408 => "00101001",
                     13409 => "00001000",
                     13410 => "11010000",
                     13411 => "00000001",
                     13412 => "11001000",
                     13413 => "10111110",
                     13414 => "01001101",
                     13415 => "10110100",
                     13416 => "10001110",
                     13417 => "00110011",
                     13418 => "00000100",
                     13419 => "10101001",
                     13420 => "00001000",
                     13421 => "10111110",
                     13422 => "01001010",
                     13423 => "10110100",
                     13424 => "10000110",
                     13425 => "10011111",
                     13426 => "00110000",
                     13427 => "00000001",
                     13428 => "01001010",
                     13429 => "10001101",
                     13430 => "00001100",
                     13431 => "00000111",
                     13432 => "01100000",
                     13433 => "10101101",
                     13434 => "00001110",
                     13435 => "00000111",
                     13436 => "11010000",
                     13437 => "00001010",
                     13438 => "10100101",
                     13439 => "00001010",
                     13440 => "00101001",
                     13441 => "10000000",
                     13442 => "11110000",
                     13443 => "00000100",
                     13444 => "00100101",
                     13445 => "00001101",
                     13446 => "11110000",
                     13447 => "00000011",
                     13448 => "01001100",
                     13449 => "00011100",
                     13450 => "10110101",
                     13451 => "10100101",
                     13452 => "00011101",
                     13453 => "11110000",
                     13454 => "00010001",
                     13455 => "10101101",
                     13456 => "00000100",
                     13457 => "00000111",
                     13458 => "11110000",
                     13459 => "11110100",
                     13460 => "10101101",
                     13461 => "10000010",
                     13462 => "00000111",
                     13463 => "11010000",
                     13464 => "00000111",
                     13465 => "10100101",
                     13466 => "10011111",
                     13467 => "00010000",
                     13468 => "00000011",
                     13469 => "01001100",
                     13470 => "00011100",
                     13471 => "10110101",
                     13472 => "10101001",
                     13473 => "00100000",
                     13474 => "10001101",
                     13475 => "10000010",
                     13476 => "00000111",
                     13477 => "10100000",
                     13478 => "00000000",
                     13479 => "10001100",
                     13480 => "00010110",
                     13481 => "00000100",
                     13482 => "10001100",
                     13483 => "00110011",
                     13484 => "00000100",
                     13485 => "10100101",
                     13486 => "10110101",
                     13487 => "10001101",
                     13488 => "00000111",
                     13489 => "00000111",
                     13490 => "10100101",
                     13491 => "11001110",
                     13492 => "10001101",
                     13493 => "00001000",
                     13494 => "00000111",
                     13495 => "10101001",
                     13496 => "00000001",
                     13497 => "10000101",
                     13498 => "00011101",
                     13499 => "10101101",
                     13500 => "00000000",
                     13501 => "00000111",
                     13502 => "11001001",
                     13503 => "00001010",
                     13504 => "10010000",
                     13505 => "00010000",
                     13506 => "11001000",
                     13507 => "11001001",
                     13508 => "00010010",
                     13509 => "10010000",
                     13510 => "00001011",
                     13511 => "11001000",
                     13512 => "11001001",
                     13513 => "00011101",
                     13514 => "10010000",
                     13515 => "00000110",
                     13516 => "11001000",
                     13517 => "11001001",
                     13518 => "00100010",
                     13519 => "10010000",
                     13520 => "00000001",
                     13521 => "11001000",
                     13522 => "10101001",
                     13523 => "00000001",
                     13524 => "10001101",
                     13525 => "00000110",
                     13526 => "00000111",
                     13527 => "10101101",
                     13528 => "00000100",
                     13529 => "00000111",
                     13530 => "11110000",
                     13531 => "00001000",
                     13532 => "10100000",
                     13533 => "00000101",
                     13534 => "10101101",
                     13535 => "01111101",
                     13536 => "00000100",
                     13537 => "11110000",
                     13538 => "00000001",
                     13539 => "11001000",
                     13540 => "10111001",
                     13541 => "00100100",
                     13542 => "10110100",
                     13543 => "10001101",
                     13544 => "00001001",
                     13545 => "00000111",
                     13546 => "10111001",
                     13547 => "00101011",
                     13548 => "10110100",
                     13549 => "10001101",
                     13550 => "00001010",
                     13551 => "00000111",
                     13552 => "10111001",
                     13553 => "00111001",
                     13554 => "10110100",
                     13555 => "10001101",
                     13556 => "00110011",
                     13557 => "00000100",
                     13558 => "10111001",
                     13559 => "00110010",
                     13560 => "10110100",
                     13561 => "10000101",
                     13562 => "10011111",
                     13563 => "10101101",
                     13564 => "00000100",
                     13565 => "00000111",
                     13566 => "11110000",
                     13567 => "00010001",
                     13568 => "10101001",
                     13569 => "00000100",
                     13570 => "10000101",
                     13571 => "11111111",
                     13572 => "10100101",
                     13573 => "11001110",
                     13574 => "11001001",
                     13575 => "00010100",
                     13576 => "10110000",
                     13577 => "00010010",
                     13578 => "10101001",
                     13579 => "00000000",
                     13580 => "10000101",
                     13581 => "10011111",
                     13582 => "01001100",
                     13583 => "00011100",
                     13584 => "10110101",
                     13585 => "10101001",
                     13586 => "00000001",
                     13587 => "10101100",
                     13588 => "01010100",
                     13589 => "00000111",
                     13590 => "11110000",
                     13591 => "00000010",
                     13592 => "10101001",
                     13593 => "10000000",
                     13594 => "10000101",
                     13595 => "11111111",
                     13596 => "10100000",
                     13597 => "00000000",
                     13598 => "10000100",
                     13599 => "00000000",
                     13600 => "10100101",
                     13601 => "00011101",
                     13602 => "11110000",
                     13603 => "00001001",
                     13604 => "10101101",
                     13605 => "00000000",
                     13606 => "00000111",
                     13607 => "11001001",
                     13608 => "00011101",
                     13609 => "10110000",
                     13610 => "00110011",
                     13611 => "10010000",
                     13612 => "00011000",
                     13613 => "11001000",
                     13614 => "10101101",
                     13615 => "01001110",
                     13616 => "00000111",
                     13617 => "11110000",
                     13618 => "00010010",
                     13619 => "10001000",
                     13620 => "10100101",
                     13621 => "00001100",
                     13622 => "11000101",
                     13623 => "01000101",
                     13624 => "11010000",
                     13625 => "00001011",
                     13626 => "10100101",
                     13627 => "00001010",
                     13628 => "00101001",
                     13629 => "01000000",
                     13630 => "11010000",
                     13631 => "00011001",
                     13632 => "10101101",
                     13633 => "10000011",
                     13634 => "00000111",
                     13635 => "11010000",
                     13636 => "00011001",
                     13637 => "11001000",
                     13638 => "11100110",
                     13639 => "00000000",
                     13640 => "10101101",
                     13641 => "00000011",
                     13642 => "00000111",
                     13643 => "11010000",
                     13644 => "00000111",
                     13645 => "10101101",
                     13646 => "00000000",
                     13647 => "00000111",
                     13648 => "11001001",
                     13649 => "00100111",
                     13650 => "10010000",
                     13651 => "00001010",
                     13652 => "11100110",
                     13653 => "00000000",
                     13654 => "01001100",
                     13655 => "01011110",
                     13656 => "10110101",
                     13657 => "10101001",
                     13658 => "00001010",
                     13659 => "10001101",
                     13660 => "10000011",
                     13661 => "00000111",
                     13662 => "10111001",
                     13663 => "01000000",
                     13664 => "10110100",
                     13665 => "10001101",
                     13666 => "01010000",
                     13667 => "00000100",
                     13668 => "10100101",
                     13669 => "00001110",
                     13670 => "11001001",
                     13671 => "00000111",
                     13672 => "11010000",
                     13673 => "00000010",
                     13674 => "10100000",
                     13675 => "00000011",
                     13676 => "10111001",
                     13677 => "01000011",
                     13678 => "10110100",
                     13679 => "10001101",
                     13680 => "01010110",
                     13681 => "00000100",
                     13682 => "10100100",
                     13683 => "00000000",
                     13684 => "10111001",
                     13685 => "01000111",
                     13686 => "10110100",
                     13687 => "10001101",
                     13688 => "00000010",
                     13689 => "00000111",
                     13690 => "10101001",
                     13691 => "00000001",
                     13692 => "10001101",
                     13693 => "00000001",
                     13694 => "00000111",
                     13695 => "10100101",
                     13696 => "00110011",
                     13697 => "11000101",
                     13698 => "01000101",
                     13699 => "11110000",
                     13700 => "00000110",
                     13701 => "00001110",
                     13702 => "00000010",
                     13703 => "00000111",
                     13704 => "00101110",
                     13705 => "00000001",
                     13706 => "00000111",
                     13707 => "01100000",
                     13708 => "00000010",
                     13709 => "00000011",
                     13710 => "00000101",
                     13711 => "10100000",
                     13712 => "00000000",
                     13713 => "10101101",
                     13714 => "00000000",
                     13715 => "00000111",
                     13716 => "11001001",
                     13717 => "00100000",
                     13718 => "10110000",
                     13719 => "00010101",
                     13720 => "11001000",
                     13721 => "11001001",
                     13722 => "00010000",
                     13723 => "10110000",
                     13724 => "00000001",
                     13725 => "11001000",
                     13726 => "10101101",
                     13727 => "11111100",
                     13728 => "00000110",
                     13729 => "00101001",
                     13730 => "01111111",
                     13731 => "11110000",
                     13732 => "00100000",
                     13733 => "00101001",
                     13734 => "00000011",
                     13735 => "11000101",
                     13736 => "01000101",
                     13737 => "11010000",
                     13738 => "00001000",
                     13739 => "10101001",
                     13740 => "00000000",
                     13741 => "10001101",
                     13742 => "00000011",
                     13743 => "00000111",
                     13744 => "01001100",
                     13745 => "11000101",
                     13746 => "10110101",
                     13747 => "10101101",
                     13748 => "00000000",
                     13749 => "00000111",
                     13750 => "11001001",
                     13751 => "00001101",
                     13752 => "10110000",
                     13753 => "00001011",
                     13754 => "10100101",
                     13755 => "00110011",
                     13756 => "10000101",
                     13757 => "01000101",
                     13758 => "10101001",
                     13759 => "00000000",
                     13760 => "10000101",
                     13761 => "01010111",
                     13762 => "10001101",
                     13763 => "00000101",
                     13764 => "00000111",
                     13765 => "10111001",
                     13766 => "10001100",
                     13767 => "10110101",
                     13768 => "10001101",
                     13769 => "00001100",
                     13770 => "00000111",
                     13771 => "01100000",
                     13772 => "00101101",
                     13773 => "10010000",
                     13774 => "00000100",
                     13775 => "11001001",
                     13776 => "00000000",
                     13777 => "11010000",
                     13778 => "00001000",
                     13779 => "10100101",
                     13780 => "01010111",
                     13781 => "11110000",
                     13782 => "01001001",
                     13783 => "00010000",
                     13784 => "00100011",
                     13785 => "00110000",
                     13786 => "00000011",
                     13787 => "01001010",
                     13788 => "10010000",
                     13789 => "00011110",
                     13790 => "10101101",
                     13791 => "00000101",
                     13792 => "00000111",
                     13793 => "00011000",
                     13794 => "01101101",
                     13795 => "00000010",
                     13796 => "00000111",
                     13797 => "10001101",
                     13798 => "00000101",
                     13799 => "00000111",
                     13800 => "10100101",
                     13801 => "01010111",
                     13802 => "01101101",
                     13803 => "00000001",
                     13804 => "00000111",
                     13805 => "10000101",
                     13806 => "01010111",
                     13807 => "11001101",
                     13808 => "01010110",
                     13809 => "00000100",
                     13810 => "00110000",
                     13811 => "00100011",
                     13812 => "10101101",
                     13813 => "01010110",
                     13814 => "00000100",
                     13815 => "10000101",
                     13816 => "01010111",
                     13817 => "01001100",
                     13818 => "00100000",
                     13819 => "10110110",
                     13820 => "10101101",
                     13821 => "00000101",
                     13822 => "00000111",
                     13823 => "00111000",
                     13824 => "11101101",
                     13825 => "00000010",
                     13826 => "00000111",
                     13827 => "10001101",
                     13828 => "00000101",
                     13829 => "00000111",
                     13830 => "10100101",
                     13831 => "01010111",
                     13832 => "11101101",
                     13833 => "00000001",
                     13834 => "00000111",
                     13835 => "10000101",
                     13836 => "01010111",
                     13837 => "11001101",
                     13838 => "01010000",
                     13839 => "00000100",
                     13840 => "00010000",
                     13841 => "00000101",
                     13842 => "10101101",
                     13843 => "01010000",
                     13844 => "00000100",
                     13845 => "10000101",
                     13846 => "01010111",
                     13847 => "11001001",
                     13848 => "00000000",
                     13849 => "00010000",
                     13850 => "00000101",
                     13851 => "01001001",
                     13852 => "11111111",
                     13853 => "00011000",
                     13854 => "01101001",
                     13855 => "00000001",
                     13856 => "10001101",
                     13857 => "00000000",
                     13858 => "00000111",
                     13859 => "01100000",
                     13860 => "10101101",
                     13861 => "01010110",
                     13862 => "00000111",
                     13863 => "11001001",
                     13864 => "00000010",
                     13865 => "10010000",
                     13866 => "01000011",
                     13867 => "10100101",
                     13868 => "00001010",
                     13869 => "00101001",
                     13870 => "01000000",
                     13871 => "11110000",
                     13872 => "00110011",
                     13873 => "00100101",
                     13874 => "00001101",
                     13875 => "11010000",
                     13876 => "00101111",
                     13877 => "10101101",
                     13878 => "11001110",
                     13879 => "00000110",
                     13880 => "00101001",
                     13881 => "00000001",
                     13882 => "10101010",
                     13883 => "10110101",
                     13884 => "00100100",
                     13885 => "11010000",
                     13886 => "00100101",
                     13887 => "10100100",
                     13888 => "10110101",
                     13889 => "10001000",
                     13890 => "11010000",
                     13891 => "00100000",
                     13892 => "10101101",
                     13893 => "00010100",
                     13894 => "00000111",
                     13895 => "11010000",
                     13896 => "00011011",
                     13897 => "10100101",
                     13898 => "00011101",
                     13899 => "11001001",
                     13900 => "00000011",
                     13901 => "11110000",
                     13902 => "00010101",
                     13903 => "10101001",
                     13904 => "00100000",
                     13905 => "10000101",
                     13906 => "11111111",
                     13907 => "10101001",
                     13908 => "00000010",
                     13909 => "10010101",
                     13910 => "00100100",
                     13911 => "10101100",
                     13912 => "00001100",
                     13913 => "00000111",
                     13914 => "10001100",
                     13915 => "00010001",
                     13916 => "00000111",
                     13917 => "10001000",
                     13918 => "10001100",
                     13919 => "10000001",
                     13920 => "00000111",
                     13921 => "11101110",
                     13922 => "11001110",
                     13923 => "00000110",
                     13924 => "10100010",
                     13925 => "00000000",
                     13926 => "00100000",
                     13927 => "10001001",
                     13928 => "10110110",
                     13929 => "10100010",
                     13930 => "00000001",
                     13931 => "00100000",
                     13932 => "10001001",
                     13933 => "10110110",
                     13934 => "10101101",
                     13935 => "01001110",
                     13936 => "00000111",
                     13937 => "11010000",
                     13938 => "00010011",
                     13939 => "10100010",
                     13940 => "00000010",
                     13941 => "10000110",
                     13942 => "00001000",
                     13943 => "00100000",
                     13944 => "11111001",
                     13945 => "10110110",
                     13946 => "00100000",
                     13947 => "00111000",
                     13948 => "11110001",
                     13949 => "00100000",
                     13950 => "10011000",
                     13951 => "11110001",
                     13952 => "00100000",
                     13953 => "11101000",
                     13954 => "11101101",
                     13955 => "11001010",
                     13956 => "00010000",
                     13957 => "11101111",
                     13958 => "01100000",
                     13959 => "01001100",
                     13960 => "10110100",
                     13961 => "10000110",
                     13962 => "00001000",
                     13963 => "10110101",
                     13964 => "00100100",
                     13965 => "00001010",
                     13966 => "10110000",
                     13967 => "01100011",
                     13968 => "10110100",
                     13969 => "00100100",
                     13970 => "11110000",
                     13971 => "01011110",
                     13972 => "10001000",
                     13973 => "11110000",
                     13974 => "00100111",
                     13975 => "10100101",
                     13976 => "10000110",
                     13977 => "01101001",
                     13978 => "00000100",
                     13979 => "10010101",
                     13980 => "10001101",
                     13981 => "10100101",
                     13982 => "01101101",
                     13983 => "01101001",
                     13984 => "00000000",
                     13985 => "10010101",
                     13986 => "01110100",
                     13987 => "10100101",
                     13988 => "11001110",
                     13989 => "10010101",
                     13990 => "11010101",
                     13991 => "10101001",
                     13992 => "00000001",
                     13993 => "10010101",
                     13994 => "10111100",
                     13995 => "10100100",
                     13996 => "00110011",
                     13997 => "10001000",
                     13998 => "10111001",
                     13999 => "10000111",
                     14000 => "10110110",
                     14001 => "10010101",
                     14002 => "01011110",
                     14003 => "10101001",
                     14004 => "00000101",
                     14005 => "10010101",
                     14006 => "10100110",
                     14007 => "10101001",
                     14008 => "00000111",
                     14009 => "10011101",
                     14010 => "10100000",
                     14011 => "00000100",
                     14012 => "11010110",
                     14013 => "00100100",
                     14014 => "10001010",
                     14015 => "00011000",
                     14016 => "01101001",
                     14017 => "00000111",
                     14018 => "10101010",
                     14019 => "10101001",
                     14020 => "01100000",
                     14021 => "10000101",
                     14022 => "00000000",
                     14023 => "10101001",
                     14024 => "00000101",
                     14025 => "10000101",
                     14026 => "00000010",
                     14027 => "10101001",
                     14028 => "00000000",
                     14029 => "00100000",
                     14030 => "11011100",
                     14031 => "10111111",
                     14032 => "00100000",
                     14033 => "00010100",
                     14034 => "10111111",
                     14035 => "10100110",
                     14036 => "00001000",
                     14037 => "00100000",
                     14038 => "01000010",
                     14039 => "11110001",
                     14040 => "00100000",
                     14041 => "10001110",
                     14042 => "11110001",
                     14043 => "00100000",
                     14044 => "00110101",
                     14045 => "11100010",
                     14046 => "00100000",
                     14047 => "11010000",
                     14048 => "11100001",
                     14049 => "10101101",
                     14050 => "11010010",
                     14051 => "00000011",
                     14052 => "00101001",
                     14053 => "11001100",
                     14054 => "11010000",
                     14055 => "00000110",
                     14056 => "00100000",
                     14057 => "11011001",
                     14058 => "11010110",
                     14059 => "01001100",
                     14060 => "11100101",
                     14061 => "11101100",
                     14062 => "10101001",
                     14063 => "00000000",
                     14064 => "10010101",
                     14065 => "00100100",
                     14066 => "01100000",
                     14067 => "00100000",
                     14068 => "01000010",
                     14069 => "11110001",
                     14070 => "01001100",
                     14071 => "00010000",
                     14072 => "11101101",
                     14073 => "10111101",
                     14074 => "10101000",
                     14075 => "00000111",
                     14076 => "00101001",
                     14077 => "00000001",
                     14078 => "10000101",
                     14079 => "00000111",
                     14080 => "10110101",
                     14081 => "11100100",
                     14082 => "11001001",
                     14083 => "11111000",
                     14084 => "11010000",
                     14085 => "00101100",
                     14086 => "10101101",
                     14087 => "10010010",
                     14088 => "00000111",
                     14089 => "11010000",
                     14090 => "00111111",
                     14091 => "10100000",
                     14092 => "00000000",
                     14093 => "10100101",
                     14094 => "00110011",
                     14095 => "01001010",
                     14096 => "10010000",
                     14097 => "00000010",
                     14098 => "10100000",
                     14099 => "00001000",
                     14100 => "10011000",
                     14101 => "01100101",
                     14102 => "10000110",
                     14103 => "10010101",
                     14104 => "10011100",
                     14105 => "10100101",
                     14106 => "01101101",
                     14107 => "01101001",
                     14108 => "00000000",
                     14109 => "10010101",
                     14110 => "10000011",
                     14111 => "10100101",
                     14112 => "11001110",
                     14113 => "00011000",
                     14114 => "01101001",
                     14115 => "00001000",
                     14116 => "10010101",
                     14117 => "11100100",
                     14118 => "10101001",
                     14119 => "00000001",
                     14120 => "10010101",
                     14121 => "11001011",
                     14122 => "10100100",
                     14123 => "00000111",
                     14124 => "10111001",
                     14125 => "01001101",
                     14126 => "10110111",
                     14127 => "10001101",
                     14128 => "10010010",
                     14129 => "00000111",
                     14130 => "10100100",
                     14131 => "00000111",
                     14132 => "10111101",
                     14133 => "00101100",
                     14134 => "00000100",
                     14135 => "00111000",
                     14136 => "11111001",
                     14137 => "01001011",
                     14138 => "10110111",
                     14139 => "10011101",
                     14140 => "00101100",
                     14141 => "00000100",
                     14142 => "10110101",
                     14143 => "11100100",
                     14144 => "11101001",
                     14145 => "00000000",
                     14146 => "11001001",
                     14147 => "00100000",
                     14148 => "10110000",
                     14149 => "00000010",
                     14150 => "10101001",
                     14151 => "11111000",
                     14152 => "10010101",
                     14153 => "11100100",
                     14154 => "01100000",
                     14155 => "11111111",
                     14156 => "01010000",
                     14157 => "01000000",
                     14158 => "00100000",
                     14159 => "10101101",
                     14160 => "01110000",
                     14161 => "00000111",
                     14162 => "11110000",
                     14163 => "01001111",
                     14164 => "10100101",
                     14165 => "00001110",
                     14166 => "11001001",
                     14167 => "00001000",
                     14168 => "10010000",
                     14169 => "01001001",
                     14170 => "11001001",
                     14171 => "00001011",
                     14172 => "11110000",
                     14173 => "01000101",
                     14174 => "10100101",
                     14175 => "10110101",
                     14176 => "11001001",
                     14177 => "00000010",
                     14178 => "10110000",
                     14179 => "00111111",
                     14180 => "10101101",
                     14181 => "10000111",
                     14182 => "00000111",
                     14183 => "11010000",
                     14184 => "00111010",
                     14185 => "10101101",
                     14186 => "11111000",
                     14187 => "00000111",
                     14188 => "00001101",
                     14189 => "11111001",
                     14190 => "00000111",
                     14191 => "00001101",
                     14192 => "11111010",
                     14193 => "00000111",
                     14194 => "11110000",
                     14195 => "00100110",
                     14196 => "10101100",
                     14197 => "11111000",
                     14198 => "00000111",
                     14199 => "10001000",
                     14200 => "11010000",
                     14201 => "00001100",
                     14202 => "10101101",
                     14203 => "11111001",
                     14204 => "00000111",
                     14205 => "00001101",
                     14206 => "11111010",
                     14207 => "00000111",
                     14208 => "11010000",
                     14209 => "00000100",
                     14210 => "10101001",
                     14211 => "01000000",
                     14212 => "10000101",
                     14213 => "11111100",
                     14214 => "10101001",
                     14215 => "00010100",
                     14216 => "10001101",
                     14217 => "10000111",
                     14218 => "00000111",
                     14219 => "10100000",
                     14220 => "00100011",
                     14221 => "10101001",
                     14222 => "11111111",
                     14223 => "10001101",
                     14224 => "00111001",
                     14225 => "00000001",
                     14226 => "00100000",
                     14227 => "01011111",
                     14228 => "10001111",
                     14229 => "10101001",
                     14230 => "10100100",
                     14231 => "01001100",
                     14232 => "00000110",
                     14233 => "10001111",
                     14234 => "10001101",
                     14235 => "01010110",
                     14236 => "00000111",
                     14237 => "00100000",
                     14238 => "00110010",
                     14239 => "11011001",
                     14240 => "11101110",
                     14241 => "01011001",
                     14242 => "00000111",
                     14243 => "01100000",
                     14244 => "10101101",
                     14245 => "00100011",
                     14246 => "00000111",
                     14247 => "11110000",
                     14248 => "11111010",
                     14249 => "10100101",
                     14250 => "11001110",
                     14251 => "00100101",
                     14252 => "10110101",
                     14253 => "11010000",
                     14254 => "11110100",
                     14255 => "10001101",
                     14256 => "00100011",
                     14257 => "00000111",
                     14258 => "11101110",
                     14259 => "11010110",
                     14260 => "00000110",
                     14261 => "01001100",
                     14262 => "10011110",
                     14263 => "11001001",
                     14264 => "10101101",
                     14265 => "01001110",
                     14266 => "00000111",
                     14267 => "11010000",
                     14268 => "00110111",
                     14269 => "10001101",
                     14270 => "01111101",
                     14271 => "00000100",
                     14272 => "10101101",
                     14273 => "01000111",
                     14274 => "00000111",
                     14275 => "11010000",
                     14276 => "00101111",
                     14277 => "10100000",
                     14278 => "00000100",
                     14279 => "10111001",
                     14280 => "01110001",
                     14281 => "00000100",
                     14282 => "00011000",
                     14283 => "01111001",
                     14284 => "01110111",
                     14285 => "00000100",
                     14286 => "10000101",
                     14287 => "00000010",
                     14288 => "10111001",
                     14289 => "01101011",
                     14290 => "00000100",
                     14291 => "11110000",
                     14292 => "00011100",
                     14293 => "01101001",
                     14294 => "00000000",
                     14295 => "10000101",
                     14296 => "00000001",
                     14297 => "10100101",
                     14298 => "10000110",
                     14299 => "00111000",
                     14300 => "11111001",
                     14301 => "01110001",
                     14302 => "00000100",
                     14303 => "10100101",
                     14304 => "01101101",
                     14305 => "11111001",
                     14306 => "01101011",
                     14307 => "00000100",
                     14308 => "00110000",
                     14309 => "00001011",
                     14310 => "10100101",
                     14311 => "00000010",
                     14312 => "00111000",
                     14313 => "11100101",
                     14314 => "10000110",
                     14315 => "10100101",
                     14316 => "00000001",
                     14317 => "11100101",
                     14318 => "01101101",
                     14319 => "00010000",
                     14320 => "00000100",
                     14321 => "10001000",
                     14322 => "00010000",
                     14323 => "11010011",
                     14324 => "01100000",
                     14325 => "10111001",
                     14326 => "01110111",
                     14327 => "00000100",
                     14328 => "01001010",
                     14329 => "10000101",
                     14330 => "00000000",
                     14331 => "10111001",
                     14332 => "01110001",
                     14333 => "00000100",
                     14334 => "00011000",
                     14335 => "01100101",
                     14336 => "00000000",
                     14337 => "10000101",
                     14338 => "00000001",
                     14339 => "10111001",
                     14340 => "01101011",
                     14341 => "00000100",
                     14342 => "01101001",
                     14343 => "00000000",
                     14344 => "10000101",
                     14345 => "00000000",
                     14346 => "10100101",
                     14347 => "00001001",
                     14348 => "01001010",
                     14349 => "10010000",
                     14350 => "00101100",
                     14351 => "10100101",
                     14352 => "00000001",
                     14353 => "00111000",
                     14354 => "11100101",
                     14355 => "10000110",
                     14356 => "10100101",
                     14357 => "00000000",
                     14358 => "11100101",
                     14359 => "01101101",
                     14360 => "00010000",
                     14361 => "00001110",
                     14362 => "10100101",
                     14363 => "10000110",
                     14364 => "00111000",
                     14365 => "11101001",
                     14366 => "00000001",
                     14367 => "10000101",
                     14368 => "10000110",
                     14369 => "10100101",
                     14370 => "01101101",
                     14371 => "11101001",
                     14372 => "00000000",
                     14373 => "01001100",
                     14374 => "00111001",
                     14375 => "10111000",
                     14376 => "10101101",
                     14377 => "10010000",
                     14378 => "00000100",
                     14379 => "01001010",
                     14380 => "10010000",
                     14381 => "00001101",
                     14382 => "10100101",
                     14383 => "10000110",
                     14384 => "00011000",
                     14385 => "01101001",
                     14386 => "00000001",
                     14387 => "10000101",
                     14388 => "10000110",
                     14389 => "10100101",
                     14390 => "01101101",
                     14391 => "01101001",
                     14392 => "00000000",
                     14393 => "10000101",
                     14394 => "01101101",
                     14395 => "10101001",
                     14396 => "00010000",
                     14397 => "10000101",
                     14398 => "00000000",
                     14399 => "10101001",
                     14400 => "00000001",
                     14401 => "10001101",
                     14402 => "01111101",
                     14403 => "00000100",
                     14404 => "10000101",
                     14405 => "00000010",
                     14406 => "01001010",
                     14407 => "10101010",
                     14408 => "01001100",
                     14409 => "11011100",
                     14410 => "10111111",
                     14411 => "00000101",
                     14412 => "00000010",
                     14413 => "00001000",
                     14414 => "00000100",
                     14415 => "00000001",
                     14416 => "00000011",
                     14417 => "00000011",
                     14418 => "00000100",
                     14419 => "00000100",
                     14420 => "00000100",
                     14421 => "10100010",
                     14422 => "00000101",
                     14423 => "10000110",
                     14424 => "00001000",
                     14425 => "10110101",
                     14426 => "00010110",
                     14427 => "11001001",
                     14428 => "00110000",
                     14429 => "11010000",
                     14430 => "01010110",
                     14431 => "10100101",
                     14432 => "00001110",
                     14433 => "11001001",
                     14434 => "00000100",
                     14435 => "11010000",
                     14436 => "00110001",
                     14437 => "10100101",
                     14438 => "00011101",
                     14439 => "11001001",
                     14440 => "00000011",
                     14441 => "11010000",
                     14442 => "00101011",
                     14443 => "10110101",
                     14444 => "11001111",
                     14445 => "11001001",
                     14446 => "10101010",
                     14447 => "10110000",
                     14448 => "00101000",
                     14449 => "10100101",
                     14450 => "11001110",
                     14451 => "11001001",
                     14452 => "10100010",
                     14453 => "10110000",
                     14454 => "00100010",
                     14455 => "10111101",
                     14456 => "00010111",
                     14457 => "00000100",
                     14458 => "01101001",
                     14459 => "11111111",
                     14460 => "10011101",
                     14461 => "00010111",
                     14462 => "00000100",
                     14463 => "10110101",
                     14464 => "11001111",
                     14465 => "01101001",
                     14466 => "00000001",
                     14467 => "10010101",
                     14468 => "11001111",
                     14469 => "10101101",
                     14470 => "00001110",
                     14471 => "00000001",
                     14472 => "00111000",
                     14473 => "11101001",
                     14474 => "11111111",
                     14475 => "10001101",
                     14476 => "00001110",
                     14477 => "00000001",
                     14478 => "10101101",
                     14479 => "00001101",
                     14480 => "00000001",
                     14481 => "11101001",
                     14482 => "00000001",
                     14483 => "10001101",
                     14484 => "00001101",
                     14485 => "00000001",
                     14486 => "01001100",
                     14487 => "10101100",
                     14488 => "10111000",
                     14489 => "10101100",
                     14490 => "00001111",
                     14491 => "00000001",
                     14492 => "10111001",
                     14493 => "01001011",
                     14494 => "10111000",
                     14495 => "10111110",
                     14496 => "01010000",
                     14497 => "10111000",
                     14498 => "10011101",
                     14499 => "00110100",
                     14500 => "00000001",
                     14501 => "00100000",
                     14502 => "00101100",
                     14503 => "10111100",
                     14504 => "10101001",
                     14505 => "00000101",
                     14506 => "10000101",
                     14507 => "00001110",
                     14508 => "00100000",
                     14509 => "10110110",
                     14510 => "11110001",
                     14511 => "00100000",
                     14512 => "01011001",
                     14513 => "11110001",
                     14514 => "00100000",
                     14515 => "01010010",
                     14516 => "11100101",
                     14517 => "01100000",
                     14518 => "00001000",
                     14519 => "00010000",
                     14520 => "00001000",
                     14521 => "00000000",
                     14522 => "00100000",
                     14523 => "10110110",
                     14524 => "11110001",
                     14525 => "10101101",
                     14526 => "01000111",
                     14527 => "00000111",
                     14528 => "11010000",
                     14529 => "01000101",
                     14530 => "10101101",
                     14531 => "00001110",
                     14532 => "00000111",
                     14533 => "11110000",
                     14534 => "01000000",
                     14535 => "10101000",
                     14536 => "10001000",
                     14537 => "10011000",
                     14538 => "00101001",
                     14539 => "00000010",
                     14540 => "11010000",
                     14541 => "00000111",
                     14542 => "11100110",
                     14543 => "11001110",
                     14544 => "11100110",
                     14545 => "11001110",
                     14546 => "01001100",
                     14547 => "11011001",
                     14548 => "10111000",
                     14549 => "11000110",
                     14550 => "11001110",
                     14551 => "11000110",
                     14552 => "11001110",
                     14553 => "10110101",
                     14554 => "01011000",
                     14555 => "00011000",
                     14556 => "01111001",
                     14557 => "10110110",
                     14558 => "10111000",
                     14559 => "10010101",
                     14560 => "11001111",
                     14561 => "11000000",
                     14562 => "00000001",
                     14563 => "10010000",
                     14564 => "00001111",
                     14565 => "10100101",
                     14566 => "00001010",
                     14567 => "00101001",
                     14568 => "10000000",
                     14569 => "11110000",
                     14570 => "00001001",
                     14571 => "00100101",
                     14572 => "00001101",
                     14573 => "11010000",
                     14574 => "00000101",
                     14575 => "10101001",
                     14576 => "11110010",
                     14577 => "10001101",
                     14578 => "11011011",
                     14579 => "00000110",
                     14580 => "11000000",
                     14581 => "00000011",
                     14582 => "11010000",
                     14583 => "00001111",
                     14584 => "10101101",
                     14585 => "11011011",
                     14586 => "00000110",
                     14587 => "10000101",
                     14588 => "10011111",
                     14589 => "10101001",
                     14590 => "01000000",
                     14591 => "10001101",
                     14592 => "00001001",
                     14593 => "00000111",
                     14594 => "10101001",
                     14595 => "00000000",
                     14596 => "10001101",
                     14597 => "00001110",
                     14598 => "00000111",
                     14599 => "00100000",
                     14600 => "01011001",
                     14601 => "11110001",
                     14602 => "00100000",
                     14603 => "10000100",
                     14604 => "11101000",
                     14605 => "00100000",
                     14606 => "01000010",
                     14607 => "11010110",
                     14608 => "10101101",
                     14609 => "00001110",
                     14610 => "00000111",
                     14611 => "11110000",
                     14612 => "00001101",
                     14613 => "10101101",
                     14614 => "10000110",
                     14615 => "00000111",
                     14616 => "11010000",
                     14617 => "00001000",
                     14618 => "10101001",
                     14619 => "00000100",
                     14620 => "10001101",
                     14621 => "10000110",
                     14622 => "00000111",
                     14623 => "11101110",
                     14624 => "00001110",
                     14625 => "00000111",
                     14626 => "01100000",
                     14627 => "10101001",
                     14628 => "00101111",
                     14629 => "10010101",
                     14630 => "00010110",
                     14631 => "10101001",
                     14632 => "00000001",
                     14633 => "10010101",
                     14634 => "00001111",
                     14635 => "10111001",
                     14636 => "01110110",
                     14637 => "00000000",
                     14638 => "10010101",
                     14639 => "01101110",
                     14640 => "10111001",
                     14641 => "10001111",
                     14642 => "00000000",
                     14643 => "10010101",
                     14644 => "10000111",
                     14645 => "10111001",
                     14646 => "11010111",
                     14647 => "00000000",
                     14648 => "10010101",
                     14649 => "11001111",
                     14650 => "10101100",
                     14651 => "10011000",
                     14652 => "00000011",
                     14653 => "11010000",
                     14654 => "00000011",
                     14655 => "10001101",
                     14656 => "10011101",
                     14657 => "00000011",
                     14658 => "10001010",
                     14659 => "10011001",
                     14660 => "10011010",
                     14661 => "00000011",
                     14662 => "11101110",
                     14663 => "10011000",
                     14664 => "00000011",
                     14665 => "10101001",
                     14666 => "00000100",
                     14667 => "10000101",
                     14668 => "11111110",
                     14669 => "01100000",
                     14670 => "00110000",
                     14671 => "01100000",
                     14672 => "11100000",
                     14673 => "00000101",
                     14674 => "11010000",
                     14675 => "01101000",
                     14676 => "10101100",
                     14677 => "10011000",
                     14678 => "00000011",
                     14679 => "10001000",
                     14680 => "10101101",
                     14681 => "10011001",
                     14682 => "00000011",
                     14683 => "11011001",
                     14684 => "01001110",
                     14685 => "10111001",
                     14686 => "11110000",
                     14687 => "00001111",
                     14688 => "10100101",
                     14689 => "00001001",
                     14690 => "01001010",
                     14691 => "01001010",
                     14692 => "10010000",
                     14693 => "00001001",
                     14694 => "10100101",
                     14695 => "11010100",
                     14696 => "11101001",
                     14697 => "00000001",
                     14698 => "10000101",
                     14699 => "11010100",
                     14700 => "11101110",
                     14701 => "10011001",
                     14702 => "00000011",
                     14703 => "10101101",
                     14704 => "10011001",
                     14705 => "00000011",
                     14706 => "11001001",
                     14707 => "00001000",
                     14708 => "10010000",
                     14709 => "01000110",
                     14710 => "00100000",
                     14711 => "01011001",
                     14712 => "11110001",
                     14713 => "00100000",
                     14714 => "10110110",
                     14715 => "11110001",
                     14716 => "10100000",
                     14717 => "00000000",
                     14718 => "00100000",
                     14719 => "00111100",
                     14720 => "11100100",
                     14721 => "11001000",
                     14722 => "11001100",
                     14723 => "10011000",
                     14724 => "00000011",
                     14725 => "11010000",
                     14726 => "11110111",
                     14727 => "10101101",
                     14728 => "11010001",
                     14729 => "00000011",
                     14730 => "00101001",
                     14731 => "00001100",
                     14732 => "11110000",
                     14733 => "00010000",
                     14734 => "10001000",
                     14735 => "10111110",
                     14736 => "10011010",
                     14737 => "00000011",
                     14738 => "00100000",
                     14739 => "10011110",
                     14740 => "11001001",
                     14741 => "10001000",
                     14742 => "00010000",
                     14743 => "11110111",
                     14744 => "10001101",
                     14745 => "10011000",
                     14746 => "00000011",
                     14747 => "10001101",
                     14748 => "10011001",
                     14749 => "00000011",
                     14750 => "10101101",
                     14751 => "10011001",
                     14752 => "00000011",
                     14753 => "11001001",
                     14754 => "00100000",
                     14755 => "10010000",
                     14756 => "00010111",
                     14757 => "10100010",
                     14758 => "00000110",
                     14759 => "10101001",
                     14760 => "00000001",
                     14761 => "10100000",
                     14762 => "00011011",
                     14763 => "00100000",
                     14764 => "11111000",
                     14765 => "11100011",
                     14766 => "10100100",
                     14767 => "00000010",
                     14768 => "11000000",
                     14769 => "11010000",
                     14770 => "10110000",
                     14771 => "00001000",
                     14772 => "10110001",
                     14773 => "00000110",
                     14774 => "11010000",
                     14775 => "00000100",
                     14776 => "10101001",
                     14777 => "00100110",
                     14778 => "10010001",
                     14779 => "00000110",
                     14780 => "10100110",
                     14781 => "00001000",
                     14782 => "01100000",
                     14783 => "00001111",
                     14784 => "00000111",
                     14785 => "10101101",
                     14786 => "01001110",
                     14787 => "00000111",
                     14788 => "11110000",
                     14789 => "01101111",
                     14790 => "10100010",
                     14791 => "00000010",
                     14792 => "10000110",
                     14793 => "00001000",
                     14794 => "10110101",
                     14795 => "00001111",
                     14796 => "11010000",
                     14797 => "01010001",
                     14798 => "10111101",
                     14799 => "10101000",
                     14800 => "00000111",
                     14801 => "10101100",
                     14802 => "11001100",
                     14803 => "00000110",
                     14804 => "00111001",
                     14805 => "10111111",
                     14806 => "10111001",
                     14807 => "11001001",
                     14808 => "00000110",
                     14809 => "10110000",
                     14810 => "01000100",
                     14811 => "10101000",
                     14812 => "10111001",
                     14813 => "01101011",
                     14814 => "00000100",
                     14815 => "11110000",
                     14816 => "00111110",
                     14817 => "10111001",
                     14818 => "01111101",
                     14819 => "00000100",
                     14820 => "11110000",
                     14821 => "00001000",
                     14822 => "11101001",
                     14823 => "00000000",
                     14824 => "10011001",
                     14825 => "01111101",
                     14826 => "00000100",
                     14827 => "01001100",
                     14828 => "00011111",
                     14829 => "10111010",
                     14830 => "10101101",
                     14831 => "01000111",
                     14832 => "00000111",
                     14833 => "11010000",
                     14834 => "00101100",
                     14835 => "10101001",
                     14836 => "00001110",
                     14837 => "10011001",
                     14838 => "01111101",
                     14839 => "00000100",
                     14840 => "10111001",
                     14841 => "01101011",
                     14842 => "00000100",
                     14843 => "10010101",
                     14844 => "01101110",
                     14845 => "10111001",
                     14846 => "01110001",
                     14847 => "00000100",
                     14848 => "10010101",
                     14849 => "10000111",
                     14850 => "10111001",
                     14851 => "01110111",
                     14852 => "00000100",
                     14853 => "00111000",
                     14854 => "11101001",
                     14855 => "00001000",
                     14856 => "10010101",
                     14857 => "11001111",
                     14858 => "10101001",
                     14859 => "00000001",
                     14860 => "10010101",
                     14861 => "10110110",
                     14862 => "10010101",
                     14863 => "00001111",
                     14864 => "01001010",
                     14865 => "10010101",
                     14866 => "00011110",
                     14867 => "10101001",
                     14868 => "00001001",
                     14869 => "10011101",
                     14870 => "10011010",
                     14871 => "00000100",
                     14872 => "10101001",
                     14873 => "00110011",
                     14874 => "10010101",
                     14875 => "00010110",
                     14876 => "01001100",
                     14877 => "00110010",
                     14878 => "10111010",
                     14879 => "10110101",
                     14880 => "00010110",
                     14881 => "11001001",
                     14882 => "00110011",
                     14883 => "11010000",
                     14884 => "00001101",
                     14885 => "00100000",
                     14886 => "01000010",
                     14887 => "11010110",
                     14888 => "10110101",
                     14889 => "00001111",
                     14890 => "11110000",
                     14891 => "00000110",
                     14892 => "00100000",
                     14893 => "10110110",
                     14894 => "11110001",
                     14895 => "00100000",
                     14896 => "00111000",
                     14897 => "10111010",
                     14898 => "11001010",
                     14899 => "00010000",
                     14900 => "10010011",
                     14901 => "01100000",
                     14902 => "00011100",
                     14903 => "11100100",
                     14904 => "10101101",
                     14905 => "01000111",
                     14906 => "00000111",
                     14907 => "11010000",
                     14908 => "00111110",
                     14909 => "10110101",
                     14910 => "00011110",
                     14911 => "11010000",
                     14912 => "00101110",
                     14913 => "10101101",
                     14914 => "11010001",
                     14915 => "00000011",
                     14916 => "00101001",
                     14917 => "00001100",
                     14918 => "11001001",
                     14919 => "00001100",
                     14920 => "11110000",
                     14921 => "01000000",
                     14922 => "10100000",
                     14923 => "00000001",
                     14924 => "00100000",
                     14925 => "01001011",
                     14926 => "11100001",
                     14927 => "00110000",
                     14928 => "00000001",
                     14929 => "11001000",
                     14930 => "10010100",
                     14931 => "01000110",
                     14932 => "10001000",
                     14933 => "10111001",
                     14934 => "00110110",
                     14935 => "10111010",
                     14936 => "10010101",
                     14937 => "01011000",
                     14938 => "10100101",
                     14939 => "00000000",
                     14940 => "01101001",
                     14941 => "00101000",
                     14942 => "11001001",
                     14943 => "01010000",
                     14944 => "10010000",
                     14945 => "00101000",
                     14946 => "10101001",
                     14947 => "00000001",
                     14948 => "10010101",
                     14949 => "00011110",
                     14950 => "10101001",
                     14951 => "00001001",
                     14952 => "10011101",
                     14953 => "10001010",
                     14954 => "00000111",
                     14955 => "10101001",
                     14956 => "00001000",
                     14957 => "10000101",
                     14958 => "11111110",
                     14959 => "10110101",
                     14960 => "00011110",
                     14961 => "00101001",
                     14962 => "00100000",
                     14963 => "11110000",
                     14964 => "00000011",
                     14965 => "00100000",
                     14966 => "01101000",
                     14967 => "10111111",
                     14968 => "00100000",
                     14969 => "00000111",
                     14970 => "10111111",
                     14971 => "00100000",
                     14972 => "10110110",
                     14973 => "11110001",
                     14974 => "00100000",
                     14975 => "01011001",
                     14976 => "11110001",
                     14977 => "00100000",
                     14978 => "01001011",
                     14979 => "11100010",
                     14980 => "00100000",
                     14981 => "01010011",
                     14982 => "11011000",
                     14983 => "01001100",
                     14984 => "10000100",
                     14985 => "11101000",
                     14986 => "00100000",
                     14987 => "10011110",
                     14988 => "11001001",
                     14989 => "01100000",
                     14990 => "00000100",
                     14991 => "00000100",
                     14992 => "00000100",
                     14993 => "00000101",
                     14994 => "00000101",
                     14995 => "00000101",
                     14996 => "00000110",
                     14997 => "00000110",
                     14998 => "00000110",
                     14999 => "00010100",
                     15000 => "11101100",
                     15001 => "10101101",
                     15002 => "10101000",
                     15003 => "00000111",
                     15004 => "00101001",
                     15005 => "00000111",
                     15006 => "11010000",
                     15007 => "00000101",
                     15008 => "10101101",
                     15009 => "10101000",
                     15010 => "00000111",
                     15011 => "00101001",
                     15012 => "00001000",
                     15013 => "10101000",
                     15014 => "10111001",
                     15015 => "00101010",
                     15016 => "00000000",
                     15017 => "11010000",
                     15018 => "00011001",
                     15019 => "10111110",
                     15020 => "10001110",
                     15021 => "10111010",
                     15022 => "10110101",
                     15023 => "00001111",
                     15024 => "11010000",
                     15025 => "00010010",
                     15026 => "10100110",
                     15027 => "00001000",
                     15028 => "10001010",
                     15029 => "10011001",
                     15030 => "10101110",
                     15031 => "00000110",
                     15032 => "10101001",
                     15033 => "10010000",
                     15034 => "10011001",
                     15035 => "00101010",
                     15036 => "00000000",
                     15037 => "10101001",
                     15038 => "00000111",
                     15039 => "10011001",
                     15040 => "10100010",
                     15041 => "00000100",
                     15042 => "00111000",
                     15043 => "01100000",
                     15044 => "10100110",
                     15045 => "00001000",
                     15046 => "00011000",
                     15047 => "01100000",
                     15048 => "10101101",
                     15049 => "01000111",
                     15050 => "00000111",
                     15051 => "11010000",
                     15052 => "01100011",
                     15053 => "10110101",
                     15054 => "00101010",
                     15055 => "00101001",
                     15056 => "01111111",
                     15057 => "10111100",
                     15058 => "10101110",
                     15059 => "00000110",
                     15060 => "11001001",
                     15061 => "00000010",
                     15062 => "11110000",
                     15063 => "00100000",
                     15064 => "10110000",
                     15065 => "00110100",
                     15066 => "10001010",
                     15067 => "00011000",
                     15068 => "01101001",
                     15069 => "00001101",
                     15070 => "10101010",
                     15071 => "10101001",
                     15072 => "00100011",
                     15073 => "10000101",
                     15074 => "00000000",
                     15075 => "10101001",
                     15076 => "00001111",
                     15077 => "10000101",
                     15078 => "00000001",
                     15079 => "10101001",
                     15080 => "00000100",
                     15081 => "10000101",
                     15082 => "00000010",
                     15083 => "10101001",
                     15084 => "00000000",
                     15085 => "00100000",
                     15086 => "11011100",
                     15087 => "10111111",
                     15088 => "00100000",
                     15089 => "00010100",
                     15090 => "10111111",
                     15091 => "10100110",
                     15092 => "00001000",
                     15093 => "01001100",
                     15094 => "00101101",
                     15095 => "10111011",
                     15096 => "10101001",
                     15097 => "11111101",
                     15098 => "10010101",
                     15099 => "10101100",
                     15100 => "10111001",
                     15101 => "00011110",
                     15102 => "00000000",
                     15103 => "00101001",
                     15104 => "11110111",
                     15105 => "10011001",
                     15106 => "00011110",
                     15107 => "00000000",
                     15108 => "10110110",
                     15109 => "01000110",
                     15110 => "11001010",
                     15111 => "10111101",
                     15112 => "10010111",
                     15113 => "10111010",
                     15114 => "10100110",
                     15115 => "00001000",
                     15116 => "10010101",
                     15117 => "01100100",
                     15118 => "11010110",
                     15119 => "00101010",
                     15120 => "10111001",
                     15121 => "10000111",
                     15122 => "00000000",
                     15123 => "00011000",
                     15124 => "01101001",
                     15125 => "00000010",
                     15126 => "10010101",
                     15127 => "10010011",
                     15128 => "10111001",
                     15129 => "01101110",
                     15130 => "00000000",
                     15131 => "01101001",
                     15132 => "00000000",
                     15133 => "10010101",
                     15134 => "01111010",
                     15135 => "10111001",
                     15136 => "11001111",
                     15137 => "00000000",
                     15138 => "00111000",
                     15139 => "11101001",
                     15140 => "00001010",
                     15141 => "10010101",
                     15142 => "11011011",
                     15143 => "10101001",
                     15144 => "00000001",
                     15145 => "10010101",
                     15146 => "11000010",
                     15147 => "11010000",
                     15148 => "00000011",
                     15149 => "00100000",
                     15150 => "11000100",
                     15151 => "11010111",
                     15152 => "00100000",
                     15153 => "10100010",
                     15154 => "11110001",
                     15155 => "00100000",
                     15156 => "01001111",
                     15157 => "11110001",
                     15158 => "00100000",
                     15159 => "00111110",
                     15160 => "11100010",
                     15161 => "00100000",
                     15162 => "11100011",
                     15163 => "11100100",
                     15164 => "01100000",
                     15165 => "00100000",
                     15166 => "10001001",
                     15167 => "10111011",
                     15168 => "10110101",
                     15169 => "01110110",
                     15170 => "10011001",
                     15171 => "01111010",
                     15172 => "00000000",
                     15173 => "10110101",
                     15174 => "10001111",
                     15175 => "00001001",
                     15176 => "00000101",
                     15177 => "10011001",
                     15178 => "10010011",
                     15179 => "00000000",
                     15180 => "10110101",
                     15181 => "11010111",
                     15182 => "11101001",
                     15183 => "00010000",
                     15184 => "10011001",
                     15185 => "11011011",
                     15186 => "00000000",
                     15187 => "01001100",
                     15188 => "01110001",
                     15189 => "10111011",
                     15190 => "00100000",
                     15191 => "10001001",
                     15192 => "10111011",
                     15193 => "10111101",
                     15194 => "11101010",
                     15195 => "00000011",
                     15196 => "10011001",
                     15197 => "01111010",
                     15198 => "00000000",
                     15199 => "10100101",
                     15200 => "00000110",
                     15201 => "00001010",
                     15202 => "00001010",
                     15203 => "00001010",
                     15204 => "00001010",
                     15205 => "00001001",
                     15206 => "00000101",
                     15207 => "10011001",
                     15208 => "10010011",
                     15209 => "00000000",
                     15210 => "10100101",
                     15211 => "00000010",
                     15212 => "01101001",
                     15213 => "00100000",
                     15214 => "10011001",
                     15215 => "11011011",
                     15216 => "00000000",
                     15217 => "10101001",
                     15218 => "11111011",
                     15219 => "10011001",
                     15220 => "10101100",
                     15221 => "00000000",
                     15222 => "10101001",
                     15223 => "00000001",
                     15224 => "10011001",
                     15225 => "11000010",
                     15226 => "00000000",
                     15227 => "10011001",
                     15228 => "00101010",
                     15229 => "00000000",
                     15230 => "10000101",
                     15231 => "11111110",
                     15232 => "10000110",
                     15233 => "00001000",
                     15234 => "00100000",
                     15235 => "00000011",
                     15236 => "10111100",
                     15237 => "11101110",
                     15238 => "01001000",
                     15239 => "00000111",
                     15240 => "01100000",
                     15241 => "10100000",
                     15242 => "00001000",
                     15243 => "10111001",
                     15244 => "00101010",
                     15245 => "00000000",
                     15246 => "11110000",
                     15247 => "00000111",
                     15248 => "10001000",
                     15249 => "11000000",
                     15250 => "00000101",
                     15251 => "11010000",
                     15252 => "11110110",
                     15253 => "10100000",
                     15254 => "00001000",
                     15255 => "10001100",
                     15256 => "10110111",
                     15257 => "00000110",
                     15258 => "01100000",
                     15259 => "10100010",
                     15260 => "00001000",
                     15261 => "10000110",
                     15262 => "00001000",
                     15263 => "10110101",
                     15264 => "00101010",
                     15265 => "11110000",
                     15266 => "01010110",
                     15267 => "00001010",
                     15268 => "10010000",
                     15269 => "00000110",
                     15270 => "00100000",
                     15271 => "11001000",
                     15272 => "10111010",
                     15273 => "01001100",
                     15274 => "11111001",
                     15275 => "10111011",
                     15276 => "10110100",
                     15277 => "00101010",
                     15278 => "10001000",
                     15279 => "11110000",
                     15280 => "00011101",
                     15281 => "11110110",
                     15282 => "00101010",
                     15283 => "10110101",
                     15284 => "10010011",
                     15285 => "00011000",
                     15286 => "01101101",
                     15287 => "01110101",
                     15288 => "00000111",
                     15289 => "10010101",
                     15290 => "10010011",
                     15291 => "10110101",
                     15292 => "01111010",
                     15293 => "01101001",
                     15294 => "00000000",
                     15295 => "10010101",
                     15296 => "01111010",
                     15297 => "10110101",
                     15298 => "00101010",
                     15299 => "11001001",
                     15300 => "00110000",
                     15301 => "11010000",
                     15302 => "00100110",
                     15303 => "10101001",
                     15304 => "00000000",
                     15305 => "10010101",
                     15306 => "00101010",
                     15307 => "01001100",
                     15308 => "11111001",
                     15309 => "10111011",
                     15310 => "10001010",
                     15311 => "00011000",
                     15312 => "01101001",
                     15313 => "00001101",
                     15314 => "10101010",
                     15315 => "10101001",
                     15316 => "01010000",
                     15317 => "10000101",
                     15318 => "00000000",
                     15319 => "10101001",
                     15320 => "00000110",
                     15321 => "10000101",
                     15322 => "00000010",
                     15323 => "01001010",
                     15324 => "10000101",
                     15325 => "00000001",
                     15326 => "10101001",
                     15327 => "00000000",
                     15328 => "00100000",
                     15329 => "11011100",
                     15330 => "10111111",
                     15331 => "10100110",
                     15332 => "00001000",
                     15333 => "10110101",
                     15334 => "10101100",
                     15335 => "11001001",
                     15336 => "00000101",
                     15337 => "11010000",
                     15338 => "00000010",
                     15339 => "11110110",
                     15340 => "00101010",
                     15341 => "00100000",
                     15342 => "01001111",
                     15343 => "11110001",
                     15344 => "00100000",
                     15345 => "10100010",
                     15346 => "11110001",
                     15347 => "00100000",
                     15348 => "00111110",
                     15349 => "11100010",
                     15350 => "00100000",
                     15351 => "10001101",
                     15352 => "11100110",
                     15353 => "11001010",
                     15354 => "00010000",
                     15355 => "10100001",
                     15356 => "01100000",
                     15357 => "00010111",
                     15358 => "00011101",
                     15359 => "00001011",
                     15360 => "00010001",
                     15361 => "00000010",
                     15362 => "00010011",
                     15363 => "10101001",
                     15364 => "00000001",
                     15365 => "10001101",
                     15366 => "00111001",
                     15367 => "00000001",
                     15368 => "10101110",
                     15369 => "01010011",
                     15370 => "00000111",
                     15371 => "10111100",
                     15372 => "11111101",
                     15373 => "10111011",
                     15374 => "00100000",
                     15375 => "01011111",
                     15376 => "10001111",
                     15377 => "11101110",
                     15378 => "01011110",
                     15379 => "00000111",
                     15380 => "10101101",
                     15381 => "01011110",
                     15382 => "00000111",
                     15383 => "11001001",
                     15384 => "01100100",
                     15385 => "11010000",
                     15386 => "00001100",
                     15387 => "10101001",
                     15388 => "00000000",
                     15389 => "10001101",
                     15390 => "01011110",
                     15391 => "00000111",
                     15392 => "11101110",
                     15393 => "01011010",
                     15394 => "00000111",
                     15395 => "10101001",
                     15396 => "01000000",
                     15397 => "10000101",
                     15398 => "11111110",
                     15399 => "10101001",
                     15400 => "00000010",
                     15401 => "10001101",
                     15402 => "00111000",
                     15403 => "00000001",
                     15404 => "10101110",
                     15405 => "01010011",
                     15406 => "00000111",
                     15407 => "10111100",
                     15408 => "11111111",
                     15409 => "10111011",
                     15410 => "00100000",
                     15411 => "01011111",
                     15412 => "10001111",
                     15413 => "10101100",
                     15414 => "01010011",
                     15415 => "00000111",
                     15416 => "10111001",
                     15417 => "00000001",
                     15418 => "10111100",
                     15419 => "00100000",
                     15420 => "00000110",
                     15421 => "10001111",
                     15422 => "10101100",
                     15423 => "00000000",
                     15424 => "00000011",
                     15425 => "10111001",
                     15426 => "11111011",
                     15427 => "00000010",
                     15428 => "11010000",
                     15429 => "00000101",
                     15430 => "10101001",
                     15431 => "00100100",
                     15432 => "10011001",
                     15433 => "11111011",
                     15434 => "00000010",
                     15435 => "10100110",
                     15436 => "00001000",
                     15437 => "01100000",
                     15438 => "10101001",
                     15439 => "00101110",
                     15440 => "10000101",
                     15441 => "00011011",
                     15442 => "10110101",
                     15443 => "01110110",
                     15444 => "10000101",
                     15445 => "01110011",
                     15446 => "10110101",
                     15447 => "10001111",
                     15448 => "10000101",
                     15449 => "10001100",
                     15450 => "10101001",
                     15451 => "00000001",
                     15452 => "10000101",
                     15453 => "10111011",
                     15454 => "10110101",
                     15455 => "11010111",
                     15456 => "00111000",
                     15457 => "11101001",
                     15458 => "00001000",
                     15459 => "10000101",
                     15460 => "11010100",
                     15461 => "10101001",
                     15462 => "00000001",
                     15463 => "10000101",
                     15464 => "00100011",
                     15465 => "10000101",
                     15466 => "00010100",
                     15467 => "10101001",
                     15468 => "00000011",
                     15469 => "10001101",
                     15470 => "10011111",
                     15471 => "00000100",
                     15472 => "10100101",
                     15473 => "00111001",
                     15474 => "11001001",
                     15475 => "00000010",
                     15476 => "10110000",
                     15477 => "00001010",
                     15478 => "10101101",
                     15479 => "01010110",
                     15480 => "00000111",
                     15481 => "11001001",
                     15482 => "00000010",
                     15483 => "10010000",
                     15484 => "00000001",
                     15485 => "01001010",
                     15486 => "10000101",
                     15487 => "00111001",
                     15488 => "10101001",
                     15489 => "00100000",
                     15490 => "10001101",
                     15491 => "11001010",
                     15492 => "00000011",
                     15493 => "10101001",
                     15494 => "00000010",
                     15495 => "10000101",
                     15496 => "11111110",
                     15497 => "01100000",
                     15498 => "10100010",
                     15499 => "00000101",
                     15500 => "10000110",
                     15501 => "00001000",
                     15502 => "10100101",
                     15503 => "00100011",
                     15504 => "11110000",
                     15505 => "01011101",
                     15506 => "00001010",
                     15507 => "10010000",
                     15508 => "00100011",
                     15509 => "10101101",
                     15510 => "01000111",
                     15511 => "00000111",
                     15512 => "11010000",
                     15513 => "01000011",
                     15514 => "10100101",
                     15515 => "00111001",
                     15516 => "11110000",
                     15517 => "00010001",
                     15518 => "11001001",
                     15519 => "00000011",
                     15520 => "11110000",
                     15521 => "00001101",
                     15522 => "11001001",
                     15523 => "00000010",
                     15524 => "11010000",
                     15525 => "00110111",
                     15526 => "00100000",
                     15527 => "11111111",
                     15528 => "11001010",
                     15529 => "00100000",
                     15530 => "01101011",
                     15531 => "11100001",
                     15532 => "01001100",
                     15533 => "11011101",
                     15534 => "10111100",
                     15535 => "00100000",
                     15536 => "01111101",
                     15537 => "11001010",
                     15538 => "00100000",
                     15539 => "11001001",
                     15540 => "11011111",
                     15541 => "01001100",
                     15542 => "11011101",
                     15543 => "10111100",
                     15544 => "10100101",
                     15545 => "00001001",
                     15546 => "00101001",
                     15547 => "00000011",
                     15548 => "11010000",
                     15549 => "00011001",
                     15550 => "11000110",
                     15551 => "11010100",
                     15552 => "10100101",
                     15553 => "00100011",
                     15554 => "11100110",
                     15555 => "00100011",
                     15556 => "11001001",
                     15557 => "00010001",
                     15558 => "10010000",
                     15559 => "00001111",
                     15560 => "10101001",
                     15561 => "00010000",
                     15562 => "10010101",
                     15563 => "01011000",
                     15564 => "10101001",
                     15565 => "10000000",
                     15566 => "10000101",
                     15567 => "00100011",
                     15568 => "00001010",
                     15569 => "10001101",
                     15570 => "11001010",
                     15571 => "00000011",
                     15572 => "00101010",
                     15573 => "10010101",
                     15574 => "01000110",
                     15575 => "10100101",
                     15576 => "00100011",
                     15577 => "11001001",
                     15578 => "00000110",
                     15579 => "10010000",
                     15580 => "00010010",
                     15581 => "00100000",
                     15582 => "01011001",
                     15583 => "11110001",
                     15584 => "00100000",
                     15585 => "10110110",
                     15586 => "11110001",
                     15587 => "00100000",
                     15588 => "01001011",
                     15589 => "11100010",
                     15590 => "00100000",
                     15591 => "11011001",
                     15592 => "11100110",
                     15593 => "00100000",
                     15594 => "01010011",
                     15595 => "11011000",
                     15596 => "00100000",
                     15597 => "01000010",
                     15598 => "11010110",
                     15599 => "01100000",
                     15600 => "00000100",
                     15601 => "00010010",
                     15602 => "01001000",
                     15603 => "10101001",
                     15604 => "00010001",
                     15605 => "10101110",
                     15606 => "11101110",
                     15607 => "00000011",
                     15608 => "10101100",
                     15609 => "01010100",
                     15610 => "00000111",
                     15611 => "11010000",
                     15612 => "00000010",
                     15613 => "10101001",
                     15614 => "00010010",
                     15615 => "10010101",
                     15616 => "00100110",
                     15617 => "00100000",
                     15618 => "01101011",
                     15619 => "10001010",
                     15620 => "10101110",
                     15621 => "11101110",
                     15622 => "00000011",
                     15623 => "10100101",
                     15624 => "00000010",
                     15625 => "10011101",
                     15626 => "11100100",
                     15627 => "00000011",
                     15628 => "10101000",
                     15629 => "10100101",
                     15630 => "00000110",
                     15631 => "10011101",
                     15632 => "11100110",
                     15633 => "00000011",
                     15634 => "10110001",
                     15635 => "00000110",
                     15636 => "00100000",
                     15637 => "11111011",
                     15638 => "10111101",
                     15639 => "10000101",
                     15640 => "00000000",
                     15641 => "10101100",
                     15642 => "01010100",
                     15643 => "00000111",
                     15644 => "11010000",
                     15645 => "00000001",
                     15646 => "10011000",
                     15647 => "10010000",
                     15648 => "00100101",
                     15649 => "10100000",
                     15650 => "00010001",
                     15651 => "10010100",
                     15652 => "00100110",
                     15653 => "10101001",
                     15654 => "11000100",
                     15655 => "10100100",
                     15656 => "00000000",
                     15657 => "11000000",
                     15658 => "01011000",
                     15659 => "11110000",
                     15660 => "00000100",
                     15661 => "11000000",
                     15662 => "01011101",
                     15663 => "11010000",
                     15664 => "00010101",
                     15665 => "10101101",
                     15666 => "10111100",
                     15667 => "00000110",
                     15668 => "11010000",
                     15669 => "00001000",
                     15670 => "10101001",
                     15671 => "00001011",
                     15672 => "10001101",
                     15673 => "10011101",
                     15674 => "00000111",
                     15675 => "11101110",
                     15676 => "10111100",
                     15677 => "00000110",
                     15678 => "10101101",
                     15679 => "10011101",
                     15680 => "00000111",
                     15681 => "11010000",
                     15682 => "00000010",
                     15683 => "10100000",
                     15684 => "11000100",
                     15685 => "10011000",
                     15686 => "10011101",
                     15687 => "11101000",
                     15688 => "00000011",
                     15689 => "00100000",
                     15690 => "10001001",
                     15691 => "10111101",
                     15692 => "10100100",
                     15693 => "00000010",
                     15694 => "10101001",
                     15695 => "00100011",
                     15696 => "10010001",
                     15697 => "00000110",
                     15698 => "10101001",
                     15699 => "00001100",
                     15700 => "10001101",
                     15701 => "10000100",
                     15702 => "00000111",
                     15703 => "01101000",
                     15704 => "10000101",
                     15705 => "00000101",
                     15706 => "10100000",
                     15707 => "00000000",
                     15708 => "10101101",
                     15709 => "00010100",
                     15710 => "00000111",
                     15711 => "11010000",
                     15712 => "00000101",
                     15713 => "10101101",
                     15714 => "01010100",
                     15715 => "00000111",
                     15716 => "11110000",
                     15717 => "00000001",
                     15718 => "11001000",
                     15719 => "10100101",
                     15720 => "11001110",
                     15721 => "00011000",
                     15722 => "01111001",
                     15723 => "11110000",
                     15724 => "10111100",
                     15725 => "00101001",
                     15726 => "11110000",
                     15727 => "10010101",
                     15728 => "11010111",
                     15729 => "10110100",
                     15730 => "00100110",
                     15731 => "11000000",
                     15732 => "00010001",
                     15733 => "11110000",
                     15734 => "00000110",
                     15735 => "00100000",
                     15736 => "00000111",
                     15737 => "10111110",
                     15738 => "01001100",
                     15739 => "10000000",
                     15740 => "10111101",
                     15741 => "00100000",
                     15742 => "10100000",
                     15743 => "10111101",
                     15744 => "10101101",
                     15745 => "11101110",
                     15746 => "00000011",
                     15747 => "01001001",
                     15748 => "00000001",
                     15749 => "10001101",
                     15750 => "11101110",
                     15751 => "00000011",
                     15752 => "01100000",
                     15753 => "10100101",
                     15754 => "10000110",
                     15755 => "00011000",
                     15756 => "01101001",
                     15757 => "00001000",
                     15758 => "00101001",
                     15759 => "11110000",
                     15760 => "10010101",
                     15761 => "10001111",
                     15762 => "10100101",
                     15763 => "01101101",
                     15764 => "01101001",
                     15765 => "00000000",
                     15766 => "10010101",
                     15767 => "01110110",
                     15768 => "10011101",
                     15769 => "11101010",
                     15770 => "00000011",
                     15771 => "10100101",
                     15772 => "10110101",
                     15773 => "10010101",
                     15774 => "10111110",
                     15775 => "01100000",
                     15776 => "00100000",
                     15777 => "00100100",
                     15778 => "10111110",
                     15779 => "10101001",
                     15780 => "00000010",
                     15781 => "10000101",
                     15782 => "11111111",
                     15783 => "10101001",
                     15784 => "00000000",
                     15785 => "10010101",
                     15786 => "01100000",
                     15787 => "10011101",
                     15788 => "00111100",
                     15789 => "00000100",
                     15790 => "10000101",
                     15791 => "10011111",
                     15792 => "10101001",
                     15793 => "11111110",
                     15794 => "10010101",
                     15795 => "10101000",
                     15796 => "10100101",
                     15797 => "00000101",
                     15798 => "00100000",
                     15799 => "11111011",
                     15800 => "10111101",
                     15801 => "10010000",
                     15802 => "00110001",
                     15803 => "10011000",
                     15804 => "11001001",
                     15805 => "00001001",
                     15806 => "10010000",
                     15807 => "00000010",
                     15808 => "11101001",
                     15809 => "00000101",
                     15810 => "00100000",
                     15811 => "00000100",
                     15812 => "10001110",
                     15813 => "11010111",
                     15814 => "10111101",
                     15815 => "00111101",
                     15816 => "10111011",
                     15817 => "00111101",
                     15818 => "10111011",
                     15819 => "11011101",
                     15820 => "10111101",
                     15821 => "11010111",
                     15822 => "10111101",
                     15823 => "11100100",
                     15824 => "10111101",
                     15825 => "11011010",
                     15826 => "10111101",
                     15827 => "00111101",
                     15828 => "10111011",
                     15829 => "11011101",
                     15830 => "10111101",
                     15831 => "10101001",
                     15832 => "00000000",
                     15833 => "00101100",
                     15834 => "10101001",
                     15835 => "00000010",
                     15836 => "00101100",
                     15837 => "10101001",
                     15838 => "00000011",
                     15839 => "10000101",
                     15840 => "00111001",
                     15841 => "01001100",
                     15842 => "01001110",
                     15843 => "10111100",
                     15844 => "10100010",
                     15845 => "00000101",
                     15846 => "10101100",
                     15847 => "11101110",
                     15848 => "00000011",
                     15849 => "00100000",
                     15850 => "00100011",
                     15851 => "10111001",
                     15852 => "01100000",
                     15853 => "11000001",
                     15854 => "11000000",
                     15855 => "01011111",
                     15856 => "01100000",
                     15857 => "01010101",
                     15858 => "01010110",
                     15859 => "01010111",
                     15860 => "01011000",
                     15861 => "01011001",
                     15862 => "01011010",
                     15863 => "01011011",
                     15864 => "01011100",
                     15865 => "01011101",
                     15866 => "01011110",
                     15867 => "10100000",
                     15868 => "00001101",
                     15869 => "11011001",
                     15870 => "11101101",
                     15871 => "10111101",
                     15872 => "11110000",
                     15873 => "00000100",
                     15874 => "10001000",
                     15875 => "00010000",
                     15876 => "11111000",
                     15877 => "00011000",
                     15878 => "01100000",
                     15879 => "00100000",
                     15880 => "00100100",
                     15881 => "10111110",
                     15882 => "10101001",
                     15883 => "00000001",
                     15884 => "10011101",
                     15885 => "11101100",
                     15886 => "00000011",
                     15887 => "10000101",
                     15888 => "11111101",
                     15889 => "00100000",
                     15890 => "01000110",
                     15891 => "10111110",
                     15892 => "10101001",
                     15893 => "11111110",
                     15894 => "10000101",
                     15895 => "10011111",
                     15896 => "10101001",
                     15897 => "00000101",
                     15898 => "10001101",
                     15899 => "00111001",
                     15900 => "00000001",
                     15901 => "00100000",
                     15902 => "00101100",
                     15903 => "10111100",
                     15904 => "10101110",
                     15905 => "11101110",
                     15906 => "00000011",
                     15907 => "01100000",
                     15908 => "10101110",
                     15909 => "11101110",
                     15910 => "00000011",
                     15911 => "10100100",
                     15912 => "00000010",
                     15913 => "11110000",
                     15914 => "00011010",
                     15915 => "10011000",
                     15916 => "00111000",
                     15917 => "11101001",
                     15918 => "00010000",
                     15919 => "10000101",
                     15920 => "00000010",
                     15921 => "10101000",
                     15922 => "10110001",
                     15923 => "00000110",
                     15924 => "11001001",
                     15925 => "11000010",
                     15926 => "11010000",
                     15927 => "00001101",
                     15928 => "10101001",
                     15929 => "00000000",
                     15930 => "10010001",
                     15931 => "00000110",
                     15932 => "00100000",
                     15933 => "01001101",
                     15934 => "10001010",
                     15935 => "10101110",
                     15936 => "11101110",
                     15937 => "00000011",
                     15938 => "00100000",
                     15939 => "01010110",
                     15940 => "10111011",
                     15941 => "01100000",
                     15942 => "10110101",
                     15943 => "10001111",
                     15944 => "10011101",
                     15945 => "11110001",
                     15946 => "00000011",
                     15947 => "10101001",
                     15948 => "11110000",
                     15949 => "10010101",
                     15950 => "01100000",
                     15951 => "10010101",
                     15952 => "01100010",
                     15953 => "10101001",
                     15954 => "11111010",
                     15955 => "10010101",
                     15956 => "10101000",
                     15957 => "10101001",
                     15958 => "11111100",
                     15959 => "10010101",
                     15960 => "10101010",
                     15961 => "10101001",
                     15962 => "00000000",
                     15963 => "10011101",
                     15964 => "00111100",
                     15965 => "00000100",
                     15966 => "10011101",
                     15967 => "00111110",
                     15968 => "00000100",
                     15969 => "10110101",
                     15970 => "01110110",
                     15971 => "10010101",
                     15972 => "01111000",
                     15973 => "10110101",
                     15974 => "10001111",
                     15975 => "10010101",
                     15976 => "10010001",
                     15977 => "10110101",
                     15978 => "11010111",
                     15979 => "00011000",
                     15980 => "01101001",
                     15981 => "00001000",
                     15982 => "10010101",
                     15983 => "11011001",
                     15984 => "10101001",
                     15985 => "11111010",
                     15986 => "10010101",
                     15987 => "10101000",
                     15988 => "01100000",
                     15989 => "10110101",
                     15990 => "00100110",
                     15991 => "11110000",
                     15992 => "01011101",
                     15993 => "00101001",
                     15994 => "00001111",
                     15995 => "01001000",
                     15996 => "10101000",
                     15997 => "10001010",
                     15998 => "00011000",
                     15999 => "01101001",
                     16000 => "00001001",
                     16001 => "10101010",
                     16002 => "10001000",
                     16003 => "11110000",
                     16004 => "00110011",
                     16005 => "00100000",
                     16006 => "10101001",
                     16007 => "10111111",
                     16008 => "00100000",
                     16009 => "00010100",
                     16010 => "10111111",
                     16011 => "10001010",
                     16012 => "00011000",
                     16013 => "01101001",
                     16014 => "00000010",
                     16015 => "10101010",
                     16016 => "00100000",
                     16017 => "10101001",
                     16018 => "10111111",
                     16019 => "00100000",
                     16020 => "00010100",
                     16021 => "10111111",
                     16022 => "10100110",
                     16023 => "00001000",
                     16024 => "00100000",
                     16025 => "01100000",
                     16026 => "11110001",
                     16027 => "00100000",
                     16028 => "10111101",
                     16029 => "11110001",
                     16030 => "00100000",
                     16031 => "01011010",
                     16032 => "11101100",
                     16033 => "01101000",
                     16034 => "10110100",
                     16035 => "10111110",
                     16036 => "11110000",
                     16037 => "00110000",
                     16038 => "01001000",
                     16039 => "10101001",
                     16040 => "11110000",
                     16041 => "11010101",
                     16042 => "11011001",
                     16043 => "10110000",
                     16044 => "00000010",
                     16045 => "10010101",
                     16046 => "11011001",
                     16047 => "10110101",
                     16048 => "11010111",
                     16049 => "11001001",
                     16050 => "11110000",
                     16051 => "01101000",
                     16052 => "10010000",
                     16053 => "00100000",
                     16054 => "10110000",
                     16055 => "00011100",
                     16056 => "00100000",
                     16057 => "10101001",
                     16058 => "10111111",
                     16059 => "10100110",
                     16060 => "00001000",
                     16061 => "00100000",
                     16062 => "01100000",
                     16063 => "11110001",
                     16064 => "00100000",
                     16065 => "10111101",
                     16066 => "11110001",
                     16067 => "00100000",
                     16068 => "11011000",
                     16069 => "11101011",
                     16070 => "10110101",
                     16071 => "11010111",
                     16072 => "00101001",
                     16073 => "00001111",
                     16074 => "11001001",
                     16075 => "00000101",
                     16076 => "01101000",
                     16077 => "10110000",
                     16078 => "00000111",
                     16079 => "10101001",
                     16080 => "00000001",
                     16081 => "10011101",
                     16082 => "11101100",
                     16083 => "00000011",
                     16084 => "10101001",
                     16085 => "00000000",
                     16086 => "10010101",
                     16087 => "00100110",
                     16088 => "01100000",
                     16089 => "10100010",
                     16090 => "00000001",
                     16091 => "10000110",
                     16092 => "00001000",
                     16093 => "10101101",
                     16094 => "00000001",
                     16095 => "00000011",
                     16096 => "11010000",
                     16097 => "00100001",
                     16098 => "10111101",
                     16099 => "11101100",
                     16100 => "00000011",
                     16101 => "11110000",
                     16102 => "00011100",
                     16103 => "10111101",
                     16104 => "11100110",
                     16105 => "00000011",
                     16106 => "10000101",
                     16107 => "00000110",
                     16108 => "10101001",
                     16109 => "00000101",
                     16110 => "10000101",
                     16111 => "00000111",
                     16112 => "10111101",
                     16113 => "11100100",
                     16114 => "00000011",
                     16115 => "10000101",
                     16116 => "00000010",
                     16117 => "10101000",
                     16118 => "10111101",
                     16119 => "11101000",
                     16120 => "00000011",
                     16121 => "10010001",
                     16122 => "00000110",
                     16123 => "00100000",
                     16124 => "01100001",
                     16125 => "10001010",
                     16126 => "10101001",
                     16127 => "00000000",
                     16128 => "10011101",
                     16129 => "11101100",
                     16130 => "00000011",
                     16131 => "11001010",
                     16132 => "00010000",
                     16133 => "11010101",
                     16134 => "01100000",
                     16135 => "11101000",
                     16136 => "00100000",
                     16137 => "00010100",
                     16138 => "10111111",
                     16139 => "10100110",
                     16140 => "00001000",
                     16141 => "01100000",
                     16142 => "10101101",
                     16143 => "00001110",
                     16144 => "00000111",
                     16145 => "11010000",
                     16146 => "00111110",
                     16147 => "10101010",
                     16148 => "10110101",
                     16149 => "01010111",
                     16150 => "00001010",
                     16151 => "00001010",
                     16152 => "00001010",
                     16153 => "00001010",
                     16154 => "10000101",
                     16155 => "00000001",
                     16156 => "10110101",
                     16157 => "01010111",
                     16158 => "01001010",
                     16159 => "01001010",
                     16160 => "01001010",
                     16161 => "01001010",
                     16162 => "11001001",
                     16163 => "00001000",
                     16164 => "10010000",
                     16165 => "00000010",
                     16166 => "00001001",
                     16167 => "11110000",
                     16168 => "10000101",
                     16169 => "00000000",
                     16170 => "10100000",
                     16171 => "00000000",
                     16172 => "11001001",
                     16173 => "00000000",
                     16174 => "00010000",
                     16175 => "00000001",
                     16176 => "10001000",
                     16177 => "10000100",
                     16178 => "00000010",
                     16179 => "10111101",
                     16180 => "00000000",
                     16181 => "00000100",
                     16182 => "00011000",
                     16183 => "01100101",
                     16184 => "00000001",
                     16185 => "10011101",
                     16186 => "00000000",
                     16187 => "00000100",
                     16188 => "10101001",
                     16189 => "00000000",
                     16190 => "00101010",
                     16191 => "01001000",
                     16192 => "01101010",
                     16193 => "10110101",
                     16194 => "10000110",
                     16195 => "01100101",
                     16196 => "00000000",
                     16197 => "10010101",
                     16198 => "10000110",
                     16199 => "10110101",
                     16200 => "01101101",
                     16201 => "01100101",
                     16202 => "00000010",
                     16203 => "10010101",
                     16204 => "01101101",
                     16205 => "01101000",
                     16206 => "00011000",
                     16207 => "01100101",
                     16208 => "00000000",
                     16209 => "01100000",
                     16210 => "10100010",
                     16211 => "00000000",
                     16212 => "10101101",
                     16213 => "01000111",
                     16214 => "00000111",
                     16215 => "11010000",
                     16216 => "00000101",
                     16217 => "10101101",
                     16218 => "00001110",
                     16219 => "00000111",
                     16220 => "11010000",
                     16221 => "11110011",
                     16222 => "10101101",
                     16223 => "00001001",
                     16224 => "00000111",
                     16225 => "10000101",
                     16226 => "00000000",
                     16227 => "10101001",
                     16228 => "00000101",
                     16229 => "01001100",
                     16230 => "10110010",
                     16231 => "10111111",
                     16232 => "10100000",
                     16233 => "00111101",
                     16234 => "10110101",
                     16235 => "00011110",
                     16236 => "11001001",
                     16237 => "00000101",
                     16238 => "11010000",
                     16239 => "00000010",
                     16240 => "10100000",
                     16241 => "00100000",
                     16242 => "01001100",
                     16243 => "10011001",
                     16244 => "10111111",
                     16245 => "10100000",
                     16246 => "00000000",
                     16247 => "01001100",
                     16248 => "01111100",
                     16249 => "10111111",
                     16250 => "10100000",
                     16251 => "00000001",
                     16252 => "11101000",
                     16253 => "10101001",
                     16254 => "00000011",
                     16255 => "10000101",
                     16256 => "00000000",
                     16257 => "10101001",
                     16258 => "00000110",
                     16259 => "10000101",
                     16260 => "00000001",
                     16261 => "10101001",
                     16262 => "00000010",
                     16263 => "10000101",
                     16264 => "00000010",
                     16265 => "10011000",
                     16266 => "01001100",
                     16267 => "11010110",
                     16268 => "10111111",
                     16269 => "10100000",
                     16270 => "01111111",
                     16271 => "11010000",
                     16272 => "00000010",
                     16273 => "10100000",
                     16274 => "00010010",
                     16275 => "10101001",
                     16276 => "00000010",
                     16277 => "11010000",
                     16278 => "00000100",
                     16279 => "10100000",
                     16280 => "00011111",
                     16281 => "10101001",
                     16282 => "00000100",
                     16283 => "10000100",
                     16284 => "00000000",
                     16285 => "11101000",
                     16286 => "00100000",
                     16287 => "10110010",
                     16288 => "10111111",
                     16289 => "10100110",
                     16290 => "00001000",
                     16291 => "01100000",
                     16292 => "00000110",
                     16293 => "00001000",
                     16294 => "10100000",
                     16295 => "00000000",
                     16296 => "00101100",
                     16297 => "10100000",
                     16298 => "00000001",
                     16299 => "10101001",
                     16300 => "01011000",
                     16301 => "10000101",
                     16302 => "00000000",
                     16303 => "10111001",
                     16304 => "10100100",
                     16305 => "10111111",
                     16306 => "10000101",
                     16307 => "00000010",
                     16308 => "10101001",
                     16309 => "00000000",
                     16310 => "01001100",
                     16311 => "11011100",
                     16312 => "10111111",
                     16313 => "10101001",
                     16314 => "00000000",
                     16315 => "00101100",
                     16316 => "10101001",
                     16317 => "00000001",
                     16318 => "01001000",
                     16319 => "10110100",
                     16320 => "00010110",
                     16321 => "11101000",
                     16322 => "10101001",
                     16323 => "00000101",
                     16324 => "11000000",
                     16325 => "00101001",
                     16326 => "11010000",
                     16327 => "00000010",
                     16328 => "10101001",
                     16329 => "00001001",
                     16330 => "10000101",
                     16331 => "00000000",
                     16332 => "10101001",
                     16333 => "00001010",
                     16334 => "10000101",
                     16335 => "00000001",
                     16336 => "10101001",
                     16337 => "00000011",
                     16338 => "10000101",
                     16339 => "00000010",
                     16340 => "01101000",
                     16341 => "10101000",
                     16342 => "00100000",
                     16343 => "11011100",
                     16344 => "10111111",
                     16345 => "10100110",
                     16346 => "00001000",
                     16347 => "01100000",
                     16348 => "01001000",
                     16349 => "10111101",
                     16350 => "00010110",
                     16351 => "00000100",
                     16352 => "00011000",
                     16353 => "01111101",
                     16354 => "00110011",
                     16355 => "00000100",
                     16356 => "10011101",
                     16357 => "00010110",
                     16358 => "00000100",
                     16359 => "10100000",
                     16360 => "00000000",
                     16361 => "10110101",
                     16362 => "10011111",
                     16363 => "00010000",
                     16364 => "00000001",
                     16365 => "10001000",
                     16366 => "10000100",
                     16367 => "00000111",
                     16368 => "01110101",
                     16369 => "11001110",
                     16370 => "10010101",
                     16371 => "11001110",
                     16372 => "10110101",
                     16373 => "10110101",
                     16374 => "01100101",
                     16375 => "00000111",
                     16376 => "10010101",
                     16377 => "10110101",
                     16378 => "10111101",
                     16379 => "00110011",
                     16380 => "00000100",
                     16381 => "00011000",
                     16382 => "01100101",
                     16383 => "00000000",
                     16384 => "10011101",
                     16385 => "00110011",
                     16386 => "00000100",
                     16387 => "10110101",
                     16388 => "10011111",
                     16389 => "01101001",
                     16390 => "00000000",
                     16391 => "10010101",
                     16392 => "10011111",
                     16393 => "11000101",
                     16394 => "00000010",
                     16395 => "00110000",
                     16396 => "00010000",
                     16397 => "10111101",
                     16398 => "00110011",
                     16399 => "00000100",
                     16400 => "11001001",
                     16401 => "10000000",
                     16402 => "10010000",
                     16403 => "00001001",
                     16404 => "10100101",
                     16405 => "00000010",
                     16406 => "10010101",
                     16407 => "10011111",
                     16408 => "10101001",
                     16409 => "00000000",
                     16410 => "10011101",
                     16411 => "00110011",
                     16412 => "00000100",
                     16413 => "01101000",
                     16414 => "11110000",
                     16415 => "00101011",
                     16416 => "10100101",
                     16417 => "00000010",
                     16418 => "01001001",
                     16419 => "11111111",
                     16420 => "10101000",
                     16421 => "11001000",
                     16422 => "10000100",
                     16423 => "00000111",
                     16424 => "10111101",
                     16425 => "00110011",
                     16426 => "00000100",
                     16427 => "00111000",
                     16428 => "11100101",
                     16429 => "00000001",
                     16430 => "10011101",
                     16431 => "00110011",
                     16432 => "00000100",
                     16433 => "10110101",
                     16434 => "10011111",
                     16435 => "11101001",
                     16436 => "00000000",
                     16437 => "10010101",
                     16438 => "10011111",
                     16439 => "11000101",
                     16440 => "00000111",
                     16441 => "00010000",
                     16442 => "00010000",
                     16443 => "10111101",
                     16444 => "00110011",
                     16445 => "00000100",
                     16446 => "11001001",
                     16447 => "10000000",
                     16448 => "10110000",
                     16449 => "00001001",
                     16450 => "10100101",
                     16451 => "00000111",
                     16452 => "10010101",
                     16453 => "10011111",
                     16454 => "10101001",
                     16455 => "11111111",
                     16456 => "10011101",
                     16457 => "00110011",
                     16458 => "00000100",
                     16459 => "01100000",
                     16460 => "11111111",
                     16461 => "10110101",
                     16462 => "00001111",
                     16463 => "01001000",
                     16464 => "00001010",
                     16465 => "10110000",
                     16466 => "00010010",
                     16467 => "01101000",
                     16468 => "11110000",
                     16469 => "00000011",
                     16470 => "01001100",
                     16471 => "10001000",
                     16472 => "11001000",
                     16473 => "10101101",
                     16474 => "00011111",
                     16475 => "00000111",
                     16476 => "00101001",
                     16477 => "00000111",
                     16478 => "11001001",
                     16479 => "00000111",
                     16480 => "11110000",
                     16481 => "00001110",
                     16482 => "01001100",
                     16483 => "11010010",
                     16484 => "11000000",
                     16485 => "01101000",
                     16486 => "00101001",
                     16487 => "00001111",
                     16488 => "10101000",
                     16489 => "10111001",
                     16490 => "00001111",
                     16491 => "00000000",
                     16492 => "11010000",
                     16493 => "00000010",
                     16494 => "10010101",
                     16495 => "00001111",
                     16496 => "01100000",
                     16497 => "00000011",
                     16498 => "00000011",
                     16499 => "00000110",
                     16500 => "00000110",
                     16501 => "00000110",
                     16502 => "00000110",
                     16503 => "00000110",
                     16504 => "00000110",
                     16505 => "00000111",
                     16506 => "00000111",
                     16507 => "00000111",
                     16508 => "00000101",
                     16509 => "00001001",
                     16510 => "00000100",
                     16511 => "00000101",
                     16512 => "00000110",
                     16513 => "00001000",
                     16514 => "00001001",
                     16515 => "00001010",
                     16516 => "00000110",
                     16517 => "00001011",
                     16518 => "00010000",
                     16519 => "01000000",
                     16520 => "10110000",
                     16521 => "10110000",
                     16522 => "10000000",
                     16523 => "01000000",
                     16524 => "01000000",
                     16525 => "10000000",
                     16526 => "01000000",
                     16527 => "11110000",
                     16528 => "11110000",
                     16529 => "11110000",
                     16530 => "10100101",
                     16531 => "01101101",
                     16532 => "00111000",
                     16533 => "11101001",
                     16534 => "00000100",
                     16535 => "10000101",
                     16536 => "01101101",
                     16537 => "10101101",
                     16538 => "00100101",
                     16539 => "00000111",
                     16540 => "00111000",
                     16541 => "11101001",
                     16542 => "00000100",
                     16543 => "10001101",
                     16544 => "00100101",
                     16545 => "00000111",
                     16546 => "10101101",
                     16547 => "00011010",
                     16548 => "00000111",
                     16549 => "00111000",
                     16550 => "11101001",
                     16551 => "00000100",
                     16552 => "10001101",
                     16553 => "00011010",
                     16554 => "00000111",
                     16555 => "10101101",
                     16556 => "00011011",
                     16557 => "00000111",
                     16558 => "00111000",
                     16559 => "11101001",
                     16560 => "00000100",
                     16561 => "10001101",
                     16562 => "00011011",
                     16563 => "00000111",
                     16564 => "10101101",
                     16565 => "00101010",
                     16566 => "00000111",
                     16567 => "00111000",
                     16568 => "11101001",
                     16569 => "00000100",
                     16570 => "10001101",
                     16571 => "00101010",
                     16572 => "00000111",
                     16573 => "10101001",
                     16574 => "00000000",
                     16575 => "10001101",
                     16576 => "00111011",
                     16577 => "00000111",
                     16578 => "10001101",
                     16579 => "00101011",
                     16580 => "00000111",
                     16581 => "10001101",
                     16582 => "00111001",
                     16583 => "00000111",
                     16584 => "10001101",
                     16585 => "00111010",
                     16586 => "00000111",
                     16587 => "10111001",
                     16588 => "11111000",
                     16589 => "10011011",
                     16590 => "10001101",
                     16591 => "00101100",
                     16592 => "00000111",
                     16593 => "01100000",
                     16594 => "10101101",
                     16595 => "01000101",
                     16596 => "00000111",
                     16597 => "11110000",
                     16598 => "01011110",
                     16599 => "10101101",
                     16600 => "00100110",
                     16601 => "00000111",
                     16602 => "11010000",
                     16603 => "01011001",
                     16604 => "10100000",
                     16605 => "00001011",
                     16606 => "10001000",
                     16607 => "00110000",
                     16608 => "01010100",
                     16609 => "10101101",
                     16610 => "01011111",
                     16611 => "00000111",
                     16612 => "11011001",
                     16613 => "01110001",
                     16614 => "11000000",
                     16615 => "11010000",
                     16616 => "11110101",
                     16617 => "10101101",
                     16618 => "00100101",
                     16619 => "00000111",
                     16620 => "11011001",
                     16621 => "01111100",
                     16622 => "11000000",
                     16623 => "11010000",
                     16624 => "11101101",
                     16625 => "10100101",
                     16626 => "11001110",
                     16627 => "11011001",
                     16628 => "10000111",
                     16629 => "11000000",
                     16630 => "11010000",
                     16631 => "00100011",
                     16632 => "10100101",
                     16633 => "00011101",
                     16634 => "11001001",
                     16635 => "00000000",
                     16636 => "11010000",
                     16637 => "00011101",
                     16638 => "10101101",
                     16639 => "01011111",
                     16640 => "00000111",
                     16641 => "11001001",
                     16642 => "00000110",
                     16643 => "11010000",
                     16644 => "00100011",
                     16645 => "11101110",
                     16646 => "11011001",
                     16647 => "00000110",
                     16648 => "11101110",
                     16649 => "11011010",
                     16650 => "00000110",
                     16651 => "10101101",
                     16652 => "11011010",
                     16653 => "00000110",
                     16654 => "11001001",
                     16655 => "00000011",
                     16656 => "11010000",
                     16657 => "00011110",
                     16658 => "10101101",
                     16659 => "11011001",
                     16660 => "00000110",
                     16661 => "11001001",
                     16662 => "00000011",
                     16663 => "11110000",
                     16664 => "00001111",
                     16665 => "11010000",
                     16666 => "00000111",
                     16667 => "10101101",
                     16668 => "01011111",
                     16669 => "00000111",
                     16670 => "11001001",
                     16671 => "00000110",
                     16672 => "11110000",
                     16673 => "11100110",
                     16674 => "00100000",
                     16675 => "10010010",
                     16676 => "11000000",
                     16677 => "00100000",
                     16678 => "00111001",
                     16679 => "11010000",
                     16680 => "10101001",
                     16681 => "00000000",
                     16682 => "10001101",
                     16683 => "11011010",
                     16684 => "00000110",
                     16685 => "10001101",
                     16686 => "11011001",
                     16687 => "00000110",
                     16688 => "10101001",
                     16689 => "00000000",
                     16690 => "10001101",
                     16691 => "01000101",
                     16692 => "00000111",
                     16693 => "10101101",
                     16694 => "11001101",
                     16695 => "00000110",
                     16696 => "11110000",
                     16697 => "00010000",
                     16698 => "10010101",
                     16699 => "00010110",
                     16700 => "10101001",
                     16701 => "00000001",
                     16702 => "10010101",
                     16703 => "00001111",
                     16704 => "10101001",
                     16705 => "00000000",
                     16706 => "10010101",
                     16707 => "00011110",
                     16708 => "10001101",
                     16709 => "11001101",
                     16710 => "00000110",
                     16711 => "01001100",
                     16712 => "00101100",
                     16713 => "11000010",
                     16714 => "10101100",
                     16715 => "00111001",
                     16716 => "00000111",
                     16717 => "10110001",
                     16718 => "11101001",
                     16719 => "11001001",
                     16720 => "11111111",
                     16721 => "11010000",
                     16722 => "00000011",
                     16723 => "01001100",
                     16724 => "00011100",
                     16725 => "11000010",
                     16726 => "00101001",
                     16727 => "00001111",
                     16728 => "11001001",
                     16729 => "00001110",
                     16730 => "11110000",
                     16731 => "00001110",
                     16732 => "11100000",
                     16733 => "00000101",
                     16734 => "10010000",
                     16735 => "00001010",
                     16736 => "11001000",
                     16737 => "10110001",
                     16738 => "11101001",
                     16739 => "00101001",
                     16740 => "00111111",
                     16741 => "11001001",
                     16742 => "00101110",
                     16743 => "11110000",
                     16744 => "00000001",
                     16745 => "01100000",
                     16746 => "10101101",
                     16747 => "00011101",
                     16748 => "00000111",
                     16749 => "00011000",
                     16750 => "01101001",
                     16751 => "00110000",
                     16752 => "00101001",
                     16753 => "11110000",
                     16754 => "10000101",
                     16755 => "00000111",
                     16756 => "10101101",
                     16757 => "00011011",
                     16758 => "00000111",
                     16759 => "01101001",
                     16760 => "00000000",
                     16761 => "10000101",
                     16762 => "00000110",
                     16763 => "10101100",
                     16764 => "00111001",
                     16765 => "00000111",
                     16766 => "11001000",
                     16767 => "10110001",
                     16768 => "11101001",
                     16769 => "00001010",
                     16770 => "10010000",
                     16771 => "00001011",
                     16772 => "10101101",
                     16773 => "00111011",
                     16774 => "00000111",
                     16775 => "11010000",
                     16776 => "00000110",
                     16777 => "11101110",
                     16778 => "00111011",
                     16779 => "00000111",
                     16780 => "11101110",
                     16781 => "00111010",
                     16782 => "00000111",
                     16783 => "10001000",
                     16784 => "10110001",
                     16785 => "11101001",
                     16786 => "00101001",
                     16787 => "00001111",
                     16788 => "11001001",
                     16789 => "00001111",
                     16790 => "11010000",
                     16791 => "00011001",
                     16792 => "10101101",
                     16793 => "00111011",
                     16794 => "00000111",
                     16795 => "11010000",
                     16796 => "00010100",
                     16797 => "11001000",
                     16798 => "10110001",
                     16799 => "11101001",
                     16800 => "00101001",
                     16801 => "00111111",
                     16802 => "10001101",
                     16803 => "00111010",
                     16804 => "00000111",
                     16805 => "11101110",
                     16806 => "00111001",
                     16807 => "00000111",
                     16808 => "11101110",
                     16809 => "00111001",
                     16810 => "00000111",
                     16811 => "11101110",
                     16812 => "00111011",
                     16813 => "00000111",
                     16814 => "01001100",
                     16815 => "11010010",
                     16816 => "11000000",
                     16817 => "10101101",
                     16818 => "00111010",
                     16819 => "00000111",
                     16820 => "10010101",
                     16821 => "01101110",
                     16822 => "10110001",
                     16823 => "11101001",
                     16824 => "00101001",
                     16825 => "11110000",
                     16826 => "10010101",
                     16827 => "10000111",
                     16828 => "11001101",
                     16829 => "00011101",
                     16830 => "00000111",
                     16831 => "10110101",
                     16832 => "01101110",
                     16833 => "11101101",
                     16834 => "00011011",
                     16835 => "00000111",
                     16836 => "10110000",
                     16837 => "00001011",
                     16838 => "10110001",
                     16839 => "11101001",
                     16840 => "00101001",
                     16841 => "00001111",
                     16842 => "11001001",
                     16843 => "00001110",
                     16844 => "11110000",
                     16845 => "01101001",
                     16846 => "01001100",
                     16847 => "01010110",
                     16848 => "11000010",
                     16849 => "10100101",
                     16850 => "00000111",
                     16851 => "11010101",
                     16852 => "10000111",
                     16853 => "10100101",
                     16854 => "00000110",
                     16855 => "11110101",
                     16856 => "01101110",
                     16857 => "10010000",
                     16858 => "01000001",
                     16859 => "10101001",
                     16860 => "00000001",
                     16861 => "10010101",
                     16862 => "10110110",
                     16863 => "10110001",
                     16864 => "11101001",
                     16865 => "00001010",
                     16866 => "00001010",
                     16867 => "00001010",
                     16868 => "00001010",
                     16869 => "10010101",
                     16870 => "11001111",
                     16871 => "11001001",
                     16872 => "11100000",
                     16873 => "11110000",
                     16874 => "01001100",
                     16875 => "11001000",
                     16876 => "10110001",
                     16877 => "11101001",
                     16878 => "00101001",
                     16879 => "01000000",
                     16880 => "11110000",
                     16881 => "00000101",
                     16882 => "10101101",
                     16883 => "11001100",
                     16884 => "00000110",
                     16885 => "11110000",
                     16886 => "01101101",
                     16887 => "10110001",
                     16888 => "11101001",
                     16889 => "00101001",
                     16890 => "00111111",
                     16891 => "11001001",
                     16892 => "00110111",
                     16893 => "10010000",
                     16894 => "00000100",
                     16895 => "11001001",
                     16896 => "00111111",
                     16897 => "10010000",
                     16898 => "00110001",
                     16899 => "11001001",
                     16900 => "00000110",
                     16901 => "11010000",
                     16902 => "00000111",
                     16903 => "10101100",
                     16904 => "01101010",
                     16905 => "00000111",
                     16906 => "11110000",
                     16907 => "00000010",
                     16908 => "10101001",
                     16909 => "00000010",
                     16910 => "10010101",
                     16911 => "00010110",
                     16912 => "10101001",
                     16913 => "00000001",
                     16914 => "10010101",
                     16915 => "00001111",
                     16916 => "00100000",
                     16917 => "00101100",
                     16918 => "11000010",
                     16919 => "10110101",
                     16920 => "00001111",
                     16921 => "11010000",
                     16922 => "01001001",
                     16923 => "01100000",
                     16924 => "10101101",
                     16925 => "11001011",
                     16926 => "00000110",
                     16927 => "11010000",
                     16928 => "00001001",
                     16929 => "10101101",
                     16930 => "10011000",
                     16931 => "00000011",
                     16932 => "11001001",
                     16933 => "00000001",
                     16934 => "11010000",
                     16935 => "00001011",
                     16936 => "10101001",
                     16937 => "00101111",
                     16938 => "10010101",
                     16939 => "00010110",
                     16940 => "10101001",
                     16941 => "00000000",
                     16942 => "10010101",
                     16943 => "00011110",
                     16944 => "00100000",
                     16945 => "01110010",
                     16946 => "11000010",
                     16947 => "01100000",
                     16948 => "01001100",
                     16949 => "00100001",
                     16950 => "11000111",
                     16951 => "11001000",
                     16952 => "11001000",
                     16953 => "10110001",
                     16954 => "11101001",
                     16955 => "01001010",
                     16956 => "01001010",
                     16957 => "01001010",
                     16958 => "01001010",
                     16959 => "01001010",
                     16960 => "11001101",
                     16961 => "01011111",
                     16962 => "00000111",
                     16963 => "11010000",
                     16964 => "00001110",
                     16965 => "10001000",
                     16966 => "10110001",
                     16967 => "11101001",
                     16968 => "10001101",
                     16969 => "01010000",
                     16970 => "00000111",
                     16971 => "11001000",
                     16972 => "10110001",
                     16973 => "11101001",
                     16974 => "00101001",
                     16975 => "00011111",
                     16976 => "10001101",
                     16977 => "01010001",
                     16978 => "00000111",
                     16979 => "01001100",
                     16980 => "01100001",
                     16981 => "11000010",
                     16982 => "10101100",
                     16983 => "00111001",
                     16984 => "00000111",
                     16985 => "10110001",
                     16986 => "11101001",
                     16987 => "00101001",
                     16988 => "00001111",
                     16989 => "11001001",
                     16990 => "00001110",
                     16991 => "11010000",
                     16992 => "00000011",
                     16993 => "11101110",
                     16994 => "00111001",
                     16995 => "00000111",
                     16996 => "11101110",
                     16997 => "00111001",
                     16998 => "00000111",
                     16999 => "11101110",
                     17000 => "00111001",
                     17001 => "00000111",
                     17002 => "10101001",
                     17003 => "00000000",
                     17004 => "10001101",
                     17005 => "00111011",
                     17006 => "00000111",
                     17007 => "10100110",
                     17008 => "00001000",
                     17009 => "01100000",
                     17010 => "10110101",
                     17011 => "00010110",
                     17012 => "11001001",
                     17013 => "00010101",
                     17014 => "10110000",
                     17015 => "00001101",
                     17016 => "10101000",
                     17017 => "10110101",
                     17018 => "11001111",
                     17019 => "01101001",
                     17020 => "00001000",
                     17021 => "10010101",
                     17022 => "11001111",
                     17023 => "10101001",
                     17024 => "00000001",
                     17025 => "10011101",
                     17026 => "11011000",
                     17027 => "00000011",
                     17028 => "10011000",
                     17029 => "00100000",
                     17030 => "00000100",
                     17031 => "10001110",
                     17032 => "00010100",
                     17033 => "11000011",
                     17034 => "00010100",
                     17035 => "11000011",
                     17036 => "00010100",
                     17037 => "11000011",
                     17038 => "00100100",
                     17039 => "11000011",
                     17040 => "11110110",
                     17041 => "11000010",
                     17042 => "00101110",
                     17043 => "11000011",
                     17044 => "11110111",
                     17045 => "11000010",
                     17046 => "01001000",
                     17047 => "11000011",
                     17048 => "01110001",
                     17049 => "11000011",
                     17050 => "11110110",
                     17051 => "11000010",
                     17052 => "01111011",
                     17053 => "11000011",
                     17054 => "01111011",
                     17055 => "11000011",
                     17056 => "11111101",
                     17057 => "11000010",
                     17058 => "10001101",
                     17059 => "11000111",
                     17060 => "11010111",
                     17061 => "11000111",
                     17062 => "01010000",
                     17063 => "11000011",
                     17064 => "01000011",
                     17065 => "11000011",
                     17066 => "10001011",
                     17067 => "11000011",
                     17068 => "10100110",
                     17069 => "11000111",
                     17070 => "11110110",
                     17071 => "11000010",
                     17072 => "10100110",
                     17073 => "11000111",
                     17074 => "10100110",
                     17075 => "11000111",
                     17076 => "10100110",
                     17077 => "11000111",
                     17078 => "10100110",
                     17079 => "11000111",
                     17080 => "10111110",
                     17081 => "11000111",
                     17082 => "11110110",
                     17083 => "11000010",
                     17084 => "11110110",
                     17085 => "11000010",
                     17086 => "01100010",
                     17087 => "11000100",
                     17088 => "01100010",
                     17089 => "11000100",
                     17090 => "01100010",
                     17091 => "11000100",
                     17092 => "01100010",
                     17093 => "11000100",
                     17094 => "01011111",
                     17095 => "11000100",
                     17096 => "11110110",
                     17097 => "11000010",
                     17098 => "11110110",
                     17099 => "11000010",
                     17100 => "11110110",
                     17101 => "11000010",
                     17102 => "11110110",
                     17103 => "11000010",
                     17104 => "11100101",
                     17105 => "11000111",
                     17106 => "00011000",
                     17107 => "11001000",
                     17108 => "01000101",
                     17109 => "11001000",
                     17110 => "01001011",
                     17111 => "11001000",
                     17112 => "00010001",
                     17113 => "11001000",
                     17114 => "00001001",
                     17115 => "11001000",
                     17116 => "00010001",
                     17117 => "11001000",
                     17118 => "01010001",
                     17119 => "11001000",
                     17120 => "01011101",
                     17121 => "11001000",
                     17122 => "01001111",
                     17123 => "11000101",
                     17124 => "01100101",
                     17125 => "10111100",
                     17126 => "00100011",
                     17127 => "10111001",
                     17128 => "11110110",
                     17129 => "11000010",
                     17130 => "11110110",
                     17131 => "11000010",
                     17132 => "11110110",
                     17133 => "11000010",
                     17134 => "11110110",
                     17135 => "11000010",
                     17136 => "11110110",
                     17137 => "11000010",
                     17138 => "00001101",
                     17139 => "11000011",
                     17140 => "10000111",
                     17141 => "11001000",
                     17142 => "01100000",
                     17143 => "00100000",
                     17144 => "00010100",
                     17145 => "11000011",
                     17146 => "01001100",
                     17147 => "01001100",
                     17148 => "11000011",
                     17149 => "10101001",
                     17150 => "00000010",
                     17151 => "10010101",
                     17152 => "10110110",
                     17153 => "10010101",
                     17154 => "11001111",
                     17155 => "01001010",
                     17156 => "10011101",
                     17157 => "10010110",
                     17158 => "00000111",
                     17159 => "01001010",
                     17160 => "10010101",
                     17161 => "00011110",
                     17162 => "01001100",
                     17163 => "01001100",
                     17164 => "11000011",
                     17165 => "10101001",
                     17166 => "10111000",
                     17167 => "10010101",
                     17168 => "11001111",
                     17169 => "01100000",
                     17170 => "11110110",
                     17171 => "11110001",
                     17172 => "10100000",
                     17173 => "00000001",
                     17174 => "10101101",
                     17175 => "01101010",
                     17176 => "00000111",
                     17177 => "11010000",
                     17178 => "00000001",
                     17179 => "10001000",
                     17180 => "10111001",
                     17181 => "00010010",
                     17182 => "11000011",
                     17183 => "10010101",
                     17184 => "01011000",
                     17185 => "01001100",
                     17186 => "01100000",
                     17187 => "11000011",
                     17188 => "00100000",
                     17189 => "00010100",
                     17190 => "11000011",
                     17191 => "10101001",
                     17192 => "00000001",
                     17193 => "10010101",
                     17194 => "00011110",
                     17195 => "01100000",
                     17196 => "10000000",
                     17197 => "01010000",
                     17198 => "10101001",
                     17199 => "00000000",
                     17200 => "10011101",
                     17201 => "10100010",
                     17202 => "00000011",
                     17203 => "10010101",
                     17204 => "01011000",
                     17205 => "10101100",
                     17206 => "11001100",
                     17207 => "00000110",
                     17208 => "10111001",
                     17209 => "00101100",
                     17210 => "11000011",
                     17211 => "10011101",
                     17212 => "10010110",
                     17213 => "00000111",
                     17214 => "10101001",
                     17215 => "00001011",
                     17216 => "01001100",
                     17217 => "01100010",
                     17218 => "11000011",
                     17219 => "10101001",
                     17220 => "00000000",
                     17221 => "01001100",
                     17222 => "00011111",
                     17223 => "11000011",
                     17224 => "10101001",
                     17225 => "00000000",
                     17226 => "10010101",
                     17227 => "01011000",
                     17228 => "10101001",
                     17229 => "00001001",
                     17230 => "11010000",
                     17231 => "00010010",
                     17232 => "10100000",
                     17233 => "00110000",
                     17234 => "10110101",
                     17235 => "11001111",
                     17236 => "10011101",
                     17237 => "00000001",
                     17238 => "00000100",
                     17239 => "00010000",
                     17240 => "00000010",
                     17241 => "10100000",
                     17242 => "11100000",
                     17243 => "10011000",
                     17244 => "01110101",
                     17245 => "11001111",
                     17246 => "10010101",
                     17247 => "01011000",
                     17248 => "10101001",
                     17249 => "00000011",
                     17250 => "10011101",
                     17251 => "10011010",
                     17252 => "00000100",
                     17253 => "10101001",
                     17254 => "00000010",
                     17255 => "10010101",
                     17256 => "01000110",
                     17257 => "10101001",
                     17258 => "00000000",
                     17259 => "10010101",
                     17260 => "10100000",
                     17261 => "10011101",
                     17262 => "00110100",
                     17263 => "00000100",
                     17264 => "01100000",
                     17265 => "10101001",
                     17266 => "00000010",
                     17267 => "10010101",
                     17268 => "01000110",
                     17269 => "10101001",
                     17270 => "00001001",
                     17271 => "10011101",
                     17272 => "10011010",
                     17273 => "00000100",
                     17274 => "01100000",
                     17275 => "00100000",
                     17276 => "01001100",
                     17277 => "11000011",
                     17278 => "10111101",
                     17279 => "10100111",
                     17280 => "00000111",
                     17281 => "00101001",
                     17282 => "00010000",
                     17283 => "10010101",
                     17284 => "01011000",
                     17285 => "10110101",
                     17286 => "11001111",
                     17287 => "10011101",
                     17288 => "00110100",
                     17289 => "00000100",
                     17290 => "01100000",
                     17291 => "10101101",
                     17292 => "11001011",
                     17293 => "00000110",
                     17294 => "11010000",
                     17295 => "00001011",
                     17296 => "10101001",
                     17297 => "00000000",
                     17298 => "10001101",
                     17299 => "11010001",
                     17300 => "00000110",
                     17301 => "00100000",
                     17302 => "01000011",
                     17303 => "11000011",
                     17304 => "01001100",
                     17305 => "11011111",
                     17306 => "11000111",
                     17307 => "01001100",
                     17308 => "10011110",
                     17309 => "11001001",
                     17310 => "00100110",
                     17311 => "00101100",
                     17312 => "00110010",
                     17313 => "00111000",
                     17314 => "00100000",
                     17315 => "00100010",
                     17316 => "00100100",
                     17317 => "00100110",
                     17318 => "00010011",
                     17319 => "00010100",
                     17320 => "00010101",
                     17321 => "00010110",
                     17322 => "10101101",
                     17323 => "10001111",
                     17324 => "00000111",
                     17325 => "11010000",
                     17326 => "00111100",
                     17327 => "11100000",
                     17328 => "00000101",
                     17329 => "10110000",
                     17330 => "00111000",
                     17331 => "10101001",
                     17332 => "10000000",
                     17333 => "10001101",
                     17334 => "10001111",
                     17335 => "00000111",
                     17336 => "10100000",
                     17337 => "00000100",
                     17338 => "10111001",
                     17339 => "00010110",
                     17340 => "00000000",
                     17341 => "11001001",
                     17342 => "00010001",
                     17343 => "11110000",
                     17344 => "00101011",
                     17345 => "10001000",
                     17346 => "00010000",
                     17347 => "11110110",
                     17348 => "11101110",
                     17349 => "11010001",
                     17350 => "00000110",
                     17351 => "10101101",
                     17352 => "11010001",
                     17353 => "00000110",
                     17354 => "11001001",
                     17355 => "00000111",
                     17356 => "10010000",
                     17357 => "00011101",
                     17358 => "10100010",
                     17359 => "00000100",
                     17360 => "10110101",
                     17361 => "00001111",
                     17362 => "11110000",
                     17363 => "00000101",
                     17364 => "11001010",
                     17365 => "00010000",
                     17366 => "11111001",
                     17367 => "00110000",
                     17368 => "00010000",
                     17369 => "10101001",
                     17370 => "00000000",
                     17371 => "10010101",
                     17372 => "00011110",
                     17373 => "10101001",
                     17374 => "00010001",
                     17375 => "10010101",
                     17376 => "00010110",
                     17377 => "00100000",
                     17378 => "10010000",
                     17379 => "11000011",
                     17380 => "10101001",
                     17381 => "00100000",
                     17382 => "00100000",
                     17383 => "11011110",
                     17384 => "11000101",
                     17385 => "10100110",
                     17386 => "00001000",
                     17387 => "01100000",
                     17388 => "10100101",
                     17389 => "11001110",
                     17390 => "11001001",
                     17391 => "00101100",
                     17392 => "10010000",
                     17393 => "11111001",
                     17394 => "10111001",
                     17395 => "00011110",
                     17396 => "00000000",
                     17397 => "11010000",
                     17398 => "11110100",
                     17399 => "10111001",
                     17400 => "01101110",
                     17401 => "00000000",
                     17402 => "10010101",
                     17403 => "01101110",
                     17404 => "10111001",
                     17405 => "10000111",
                     17406 => "00000000",
                     17407 => "10010101",
                     17408 => "10000111",
                     17409 => "10101001",
                     17410 => "00000001",
                     17411 => "10010101",
                     17412 => "10110110",
                     17413 => "10111001",
                     17414 => "11001111",
                     17415 => "00000000",
                     17416 => "00111000",
                     17417 => "11101001",
                     17418 => "00001000",
                     17419 => "10010101",
                     17420 => "11001111",
                     17421 => "10111101",
                     17422 => "10100111",
                     17423 => "00000111",
                     17424 => "00101001",
                     17425 => "00000011",
                     17426 => "10101000",
                     17427 => "10100010",
                     17428 => "00000010",
                     17429 => "10111001",
                     17430 => "10011110",
                     17431 => "11000011",
                     17432 => "10010101",
                     17433 => "00000001",
                     17434 => "11001000",
                     17435 => "11001000",
                     17436 => "11001000",
                     17437 => "11001000",
                     17438 => "11001010",
                     17439 => "00010000",
                     17440 => "11110100",
                     17441 => "10100110",
                     17442 => "00001000",
                     17443 => "00100000",
                     17444 => "00110100",
                     17445 => "11001111",
                     17446 => "10100100",
                     17447 => "01010111",
                     17448 => "11000000",
                     17449 => "00001100",
                     17450 => "10110000",
                     17451 => "00001110",
                     17452 => "10101000",
                     17453 => "10111101",
                     17454 => "10101000",
                     17455 => "00000111",
                     17456 => "00101001",
                     17457 => "00000011",
                     17458 => "11110000",
                     17459 => "00000101",
                     17460 => "10011000",
                     17461 => "01001001",
                     17462 => "11111111",
                     17463 => "10101000",
                     17464 => "11001000",
                     17465 => "10011000",
                     17466 => "00100000",
                     17467 => "01001100",
                     17468 => "11000011",
                     17469 => "10100000",
                     17470 => "00000010",
                     17471 => "10010101",
                     17472 => "01011000",
                     17473 => "11001001",
                     17474 => "00000000",
                     17475 => "00110000",
                     17476 => "00000001",
                     17477 => "10001000",
                     17478 => "10010100",
                     17479 => "01000110",
                     17480 => "10101001",
                     17481 => "11111101",
                     17482 => "10010101",
                     17483 => "10100000",
                     17484 => "10101001",
                     17485 => "00000001",
                     17486 => "10010101",
                     17487 => "00001111",
                     17488 => "10101001",
                     17489 => "00000101",
                     17490 => "10010101",
                     17491 => "00011110",
                     17492 => "01100000",
                     17493 => "00110000",
                     17494 => "01000011",
                     17495 => "00110000",
                     17496 => "01000011",
                     17497 => "00110000",
                     17498 => "00000000",
                     17499 => "00000000",
                     17500 => "00010000",
                     17501 => "00010000",
                     17502 => "00000000",
                     17503 => "00100000",
                     17504 => "01111011",
                     17505 => "11000101",
                     17506 => "10101001",
                     17507 => "00000000",
                     17508 => "10010101",
                     17509 => "01011000",
                     17510 => "10110101",
                     17511 => "00010110",
                     17512 => "00111000",
                     17513 => "11101001",
                     17514 => "00011011",
                     17515 => "10101000",
                     17516 => "10111001",
                     17517 => "01010101",
                     17518 => "11000100",
                     17519 => "10011101",
                     17520 => "10001000",
                     17521 => "00000011",
                     17522 => "10111001",
                     17523 => "01011010",
                     17524 => "11000100",
                     17525 => "10010101",
                     17526 => "00110100",
                     17527 => "10110101",
                     17528 => "11001111",
                     17529 => "00011000",
                     17530 => "01101001",
                     17531 => "00000100",
                     17532 => "10010101",
                     17533 => "11001111",
                     17534 => "10110101",
                     17535 => "10000111",
                     17536 => "00011000",
                     17537 => "01101001",
                     17538 => "00000100",
                     17539 => "10010101",
                     17540 => "10000111",
                     17541 => "10110101",
                     17542 => "01101110",
                     17543 => "01101001",
                     17544 => "00000000",
                     17545 => "10010101",
                     17546 => "01101110",
                     17547 => "01001100",
                     17548 => "11011111",
                     17549 => "11000111",
                     17550 => "10000000",
                     17551 => "00110000",
                     17552 => "01000000",
                     17553 => "10000000",
                     17554 => "00110000",
                     17555 => "01010000",
                     17556 => "01010000",
                     17557 => "01110000",
                     17558 => "00100000",
                     17559 => "01000000",
                     17560 => "10000000",
                     17561 => "10100000",
                     17562 => "01110000",
                     17563 => "01000000",
                     17564 => "10010000",
                     17565 => "01101000",
                     17566 => "00010001",
                     17567 => "00000111",
                     17568 => "00001000",
                     17569 => "00001010",
                     17570 => "00100011",
                     17571 => "00101000",
                     17572 => "00010101",
                     17573 => "00010000",
                     17574 => "00100010",
                     17575 => "00101100",
                     17576 => "00011111",
                     17577 => "00011011",
                     17578 => "00010000",
                     17579 => "01100000",
                     17580 => "00100000",
                     17581 => "01001000",
                     17582 => "10101101",
                     17583 => "10001111",
                     17584 => "00000111",
                     17585 => "11010000",
                     17586 => "10100001",
                     17587 => "00100000",
                     17588 => "01001100",
                     17589 => "11000011",
                     17590 => "10111101",
                     17591 => "10101000",
                     17592 => "00000111",
                     17593 => "00101001",
                     17594 => "00000011",
                     17595 => "10101000",
                     17596 => "10111001",
                     17597 => "10101010",
                     17598 => "11000100",
                     17599 => "10001101",
                     17600 => "10001111",
                     17601 => "00000111",
                     17602 => "10100000",
                     17603 => "00000011",
                     17604 => "10101101",
                     17605 => "11001100",
                     17606 => "00000110",
                     17607 => "11110000",
                     17608 => "00000001",
                     17609 => "11001000",
                     17610 => "10000100",
                     17611 => "00000000",
                     17612 => "11100100",
                     17613 => "00000000",
                     17614 => "10110000",
                     17615 => "10000100",
                     17616 => "10111101",
                     17617 => "10100111",
                     17618 => "00000111",
                     17619 => "00101001",
                     17620 => "00000011",
                     17621 => "10000101",
                     17622 => "00000000",
                     17623 => "10000101",
                     17624 => "00000001",
                     17625 => "10101001",
                     17626 => "11111010",
                     17627 => "10010101",
                     17628 => "10100000",
                     17629 => "10101001",
                     17630 => "00000000",
                     17631 => "10100100",
                     17632 => "01010111",
                     17633 => "11110000",
                     17634 => "00000111",
                     17635 => "10101001",
                     17636 => "00000100",
                     17637 => "11000000",
                     17638 => "00011101",
                     17639 => "10010000",
                     17640 => "00000001",
                     17641 => "00001010",
                     17642 => "01001000",
                     17643 => "00011000",
                     17644 => "01100101",
                     17645 => "00000000",
                     17646 => "10000101",
                     17647 => "00000000",
                     17648 => "10111101",
                     17649 => "10101000",
                     17650 => "00000111",
                     17651 => "00101001",
                     17652 => "00000011",
                     17653 => "11110000",
                     17654 => "00000111",
                     17655 => "10111101",
                     17656 => "10101001",
                     17657 => "00000111",
                     17658 => "00101001",
                     17659 => "00001111",
                     17660 => "10000101",
                     17661 => "00000000",
                     17662 => "01101000",
                     17663 => "00011000",
                     17664 => "01100101",
                     17665 => "00000001",
                     17666 => "10101000",
                     17667 => "10111001",
                     17668 => "10011110",
                     17669 => "11000100",
                     17670 => "10010101",
                     17671 => "01011000",
                     17672 => "10101001",
                     17673 => "00000001",
                     17674 => "10010101",
                     17675 => "01000110",
                     17676 => "10100101",
                     17677 => "01010111",
                     17678 => "11010000",
                     17679 => "00010010",
                     17680 => "10100100",
                     17681 => "00000000",
                     17682 => "10011000",
                     17683 => "00101001",
                     17684 => "00000010",
                     17685 => "11110000",
                     17686 => "00001011",
                     17687 => "10110101",
                     17688 => "01011000",
                     17689 => "01001001",
                     17690 => "11111111",
                     17691 => "00011000",
                     17692 => "01101001",
                     17693 => "00000001",
                     17694 => "10010101",
                     17695 => "01011000",
                     17696 => "11110110",
                     17697 => "01000110",
                     17698 => "10011000",
                     17699 => "00101001",
                     17700 => "00000010",
                     17701 => "11110000",
                     17702 => "00001111",
                     17703 => "10100101",
                     17704 => "10000110",
                     17705 => "00011000",
                     17706 => "01111001",
                     17707 => "10001110",
                     17708 => "11000100",
                     17709 => "10010101",
                     17710 => "10000111",
                     17711 => "10100101",
                     17712 => "01101101",
                     17713 => "01101001",
                     17714 => "00000000",
                     17715 => "01001100",
                     17716 => "01000010",
                     17717 => "11000101",
                     17718 => "10100101",
                     17719 => "10000110",
                     17720 => "00111000",
                     17721 => "11111001",
                     17722 => "10001110",
                     17723 => "11000100",
                     17724 => "10010101",
                     17725 => "10000111",
                     17726 => "10100101",
                     17727 => "01101101",
                     17728 => "11101001",
                     17729 => "00000000",
                     17730 => "10010101",
                     17731 => "01101110",
                     17732 => "10101001",
                     17733 => "00000001",
                     17734 => "10010101",
                     17735 => "00001111",
                     17736 => "10010101",
                     17737 => "10110110",
                     17738 => "10101001",
                     17739 => "11111000",
                     17740 => "10010101",
                     17741 => "11001111",
                     17742 => "01100000",
                     17743 => "00100000",
                     17744 => "01111011",
                     17745 => "11000101",
                     17746 => "10001110",
                     17747 => "01101000",
                     17748 => "00000011",
                     17749 => "10101001",
                     17750 => "00000000",
                     17751 => "10001101",
                     17752 => "01100011",
                     17753 => "00000011",
                     17754 => "10001101",
                     17755 => "01101001",
                     17756 => "00000011",
                     17757 => "10110101",
                     17758 => "10000111",
                     17759 => "10001101",
                     17760 => "01100110",
                     17761 => "00000011",
                     17762 => "10101001",
                     17763 => "11011111",
                     17764 => "10001101",
                     17765 => "10010000",
                     17766 => "00000111",
                     17767 => "10010101",
                     17768 => "01000110",
                     17769 => "10101001",
                     17770 => "00100000",
                     17771 => "10001101",
                     17772 => "01100100",
                     17773 => "00000011",
                     17774 => "10011101",
                     17775 => "10001010",
                     17776 => "00000111",
                     17777 => "10101001",
                     17778 => "00000101",
                     17779 => "10001101",
                     17780 => "10000011",
                     17781 => "00000100",
                     17782 => "01001010",
                     17783 => "10001101",
                     17784 => "01100101",
                     17785 => "00000011",
                     17786 => "01100000",
                     17787 => "10100000",
                     17788 => "11111111",
                     17789 => "11001000",
                     17790 => "10111001",
                     17791 => "00001111",
                     17792 => "00000000",
                     17793 => "11010000",
                     17794 => "11111010",
                     17795 => "10001100",
                     17796 => "11001111",
                     17797 => "00000110",
                     17798 => "10001010",
                     17799 => "00001001",
                     17800 => "10000000",
                     17801 => "10011001",
                     17802 => "00001111",
                     17803 => "00000000",
                     17804 => "10110101",
                     17805 => "01101110",
                     17806 => "10011001",
                     17807 => "01101110",
                     17808 => "00000000",
                     17809 => "10110101",
                     17810 => "10000111",
                     17811 => "10011001",
                     17812 => "10000111",
                     17813 => "00000000",
                     17814 => "10101001",
                     17815 => "00000001",
                     17816 => "10010101",
                     17817 => "00001111",
                     17818 => "10011001",
                     17819 => "10110110",
                     17820 => "00000000",
                     17821 => "10110101",
                     17822 => "11001111",
                     17823 => "10011001",
                     17824 => "11001111",
                     17825 => "00000000",
                     17826 => "01100000",
                     17827 => "10010000",
                     17828 => "10000000",
                     17829 => "01110000",
                     17830 => "10010000",
                     17831 => "11111111",
                     17832 => "00000001",
                     17833 => "10101101",
                     17834 => "10001111",
                     17835 => "00000111",
                     17836 => "11010000",
                     17837 => "11110100",
                     17838 => "10011101",
                     17839 => "00110100",
                     17840 => "00000100",
                     17841 => "10100101",
                     17842 => "11111101",
                     17843 => "00001001",
                     17844 => "00000010",
                     17845 => "10000101",
                     17846 => "11111101",
                     17847 => "10101100",
                     17848 => "01101000",
                     17849 => "00000011",
                     17850 => "10111001",
                     17851 => "00010110",
                     17852 => "00000000",
                     17853 => "11001001",
                     17854 => "00101101",
                     17855 => "11110000",
                     17856 => "00110001",
                     17857 => "00100000",
                     17858 => "10100001",
                     17859 => "11010001",
                     17860 => "00011000",
                     17861 => "01101001",
                     17862 => "00100000",
                     17863 => "10101100",
                     17864 => "11001100",
                     17865 => "00000110",
                     17866 => "11110000",
                     17867 => "00000011",
                     17868 => "00111000",
                     17869 => "11101001",
                     17870 => "00010000",
                     17871 => "10001101",
                     17872 => "10001111",
                     17873 => "00000111",
                     17874 => "10111101",
                     17875 => "10100111",
                     17876 => "00000111",
                     17877 => "00101001",
                     17878 => "00000011",
                     17879 => "10011101",
                     17880 => "00010111",
                     17881 => "00000100",
                     17882 => "10101000",
                     17883 => "10111001",
                     17884 => "10100011",
                     17885 => "11000101",
                     17886 => "10010101",
                     17887 => "11001111",
                     17888 => "10101101",
                     17889 => "00011101",
                     17890 => "00000111",
                     17891 => "00011000",
                     17892 => "01101001",
                     17893 => "00100000",
                     17894 => "10010101",
                     17895 => "10000111",
                     17896 => "10101101",
                     17897 => "00011011",
                     17898 => "00000111",
                     17899 => "01101001",
                     17900 => "00000000",
                     17901 => "10010101",
                     17902 => "01101110",
                     17903 => "01001100",
                     17904 => "00100101",
                     17905 => "11000110",
                     17906 => "10111001",
                     17907 => "10000111",
                     17908 => "00000000",
                     17909 => "00111000",
                     17910 => "11101001",
                     17911 => "00001110",
                     17912 => "10010101",
                     17913 => "10000111",
                     17914 => "10111001",
                     17915 => "01101110",
                     17916 => "00000000",
                     17917 => "10010101",
                     17918 => "01101110",
                     17919 => "10111001",
                     17920 => "11001111",
                     17921 => "00000000",
                     17922 => "00011000",
                     17923 => "01101001",
                     17924 => "00001000",
                     17925 => "10010101",
                     17926 => "11001111",
                     17927 => "10111101",
                     17928 => "10100111",
                     17929 => "00000111",
                     17930 => "00101001",
                     17931 => "00000011",
                     17932 => "10011101",
                     17933 => "00010111",
                     17934 => "00000100",
                     17935 => "10101000",
                     17936 => "10111001",
                     17937 => "10100011",
                     17938 => "11000101",
                     17939 => "10100000",
                     17940 => "00000000",
                     17941 => "11010101",
                     17942 => "11001111",
                     17943 => "10010000",
                     17944 => "00000001",
                     17945 => "11001000",
                     17946 => "10111001",
                     17947 => "10100111",
                     17948 => "11000101",
                     17949 => "10011101",
                     17950 => "00110100",
                     17951 => "00000100",
                     17952 => "10101001",
                     17953 => "00000000",
                     17954 => "10001101",
                     17955 => "11001011",
                     17956 => "00000110",
                     17957 => "10101001",
                     17958 => "00001000",
                     17959 => "10011101",
                     17960 => "10011010",
                     17961 => "00000100",
                     17962 => "10101001",
                     17963 => "00000001",
                     17964 => "10010101",
                     17965 => "10110110",
                     17966 => "10010101",
                     17967 => "00001111",
                     17968 => "01001010",
                     17969 => "10011101",
                     17970 => "00000001",
                     17971 => "00000100",
                     17972 => "10010101",
                     17973 => "00011110",
                     17974 => "01100000",
                     17975 => "00000000",
                     17976 => "00110000",
                     17977 => "01100000",
                     17978 => "01100000",
                     17979 => "00000000",
                     17980 => "00100000",
                     17981 => "01100000",
                     17982 => "01000000",
                     17983 => "01110000",
                     17984 => "01000000",
                     17985 => "01100000",
                     17986 => "00110000",
                     17987 => "10101101",
                     17988 => "10001111",
                     17989 => "00000111",
                     17990 => "11010000",
                     17991 => "01000111",
                     17992 => "10101001",
                     17993 => "00100000",
                     17994 => "10001101",
                     17995 => "10001111",
                     17996 => "00000111",
                     17997 => "11001110",
                     17998 => "11010111",
                     17999 => "00000110",
                     18000 => "10100000",
                     18001 => "00000110",
                     18002 => "10001000",
                     18003 => "10111001",
                     18004 => "00010110",
                     18005 => "00000000",
                     18006 => "11001001",
                     18007 => "00110001",
                     18008 => "11010000",
                     18009 => "11111000",
                     18010 => "10111001",
                     18011 => "10000111",
                     18012 => "00000000",
                     18013 => "00111000",
                     18014 => "11101001",
                     18015 => "00110000",
                     18016 => "01001000",
                     18017 => "10111001",
                     18018 => "01101110",
                     18019 => "00000000",
                     18020 => "11101001",
                     18021 => "00000000",
                     18022 => "10000101",
                     18023 => "00000000",
                     18024 => "10101101",
                     18025 => "11010111",
                     18026 => "00000110",
                     18027 => "00011000",
                     18028 => "01111001",
                     18029 => "00011110",
                     18030 => "00000000",
                     18031 => "10101000",
                     18032 => "01101000",
                     18033 => "00011000",
                     18034 => "01111001",
                     18035 => "00110111",
                     18036 => "11000110",
                     18037 => "10010101",
                     18038 => "10000111",
                     18039 => "10100101",
                     18040 => "00000000",
                     18041 => "01101001",
                     18042 => "00000000",
                     18043 => "10010101",
                     18044 => "01101110",
                     18045 => "10111001",
                     18046 => "00111101",
                     18047 => "11000110",
                     18048 => "10010101",
                     18049 => "11001111",
                     18050 => "10101001",
                     18051 => "00000001",
                     18052 => "10010101",
                     18053 => "10110110",
                     18054 => "10010101",
                     18055 => "00001111",
                     18056 => "01001010",
                     18057 => "10010101",
                     18058 => "01011000",
                     18059 => "10101001",
                     18060 => "00001000",
                     18061 => "10010101",
                     18062 => "10100000",
                     18063 => "01100000",
                     18064 => "00000001",
                     18065 => "00000010",
                     18066 => "00000100",
                     18067 => "00001000",
                     18068 => "00010000",
                     18069 => "00100000",
                     18070 => "01000000",
                     18071 => "10000000",
                     18072 => "01000000",
                     18073 => "00110000",
                     18074 => "10010000",
                     18075 => "01010000",
                     18076 => "00100000",
                     18077 => "01100000",
                     18078 => "10100000",
                     18079 => "01110000",
                     18080 => "00001010",
                     18081 => "00001011",
                     18082 => "10101101",
                     18083 => "10001111",
                     18084 => "00000111",
                     18085 => "11010000",
                     18086 => "01101111",
                     18087 => "10101101",
                     18088 => "01001110",
                     18089 => "00000111",
                     18090 => "11010000",
                     18091 => "01010111",
                     18092 => "11100000",
                     18093 => "00000011",
                     18094 => "10110000",
                     18095 => "01100110",
                     18096 => "10100000",
                     18097 => "00000000",
                     18098 => "10111101",
                     18099 => "10100111",
                     18100 => "00000111",
                     18101 => "11001001",
                     18102 => "10101010",
                     18103 => "10010000",
                     18104 => "00000001",
                     18105 => "11001000",
                     18106 => "10101101",
                     18107 => "01011111",
                     18108 => "00000111",
                     18109 => "11001001",
                     18110 => "00000001",
                     18111 => "11110000",
                     18112 => "00000001",
                     18113 => "11001000",
                     18114 => "10011000",
                     18115 => "00101001",
                     18116 => "00000001",
                     18117 => "10101000",
                     18118 => "10111001",
                     18119 => "10100000",
                     18120 => "11000110",
                     18121 => "10010101",
                     18122 => "00010110",
                     18123 => "10101101",
                     18124 => "11011101",
                     18125 => "00000110",
                     18126 => "11001001",
                     18127 => "11111111",
                     18128 => "11010000",
                     18129 => "00000101",
                     18130 => "10101001",
                     18131 => "00000000",
                     18132 => "10001101",
                     18133 => "11011101",
                     18134 => "00000110",
                     18135 => "10111101",
                     18136 => "10100111",
                     18137 => "00000111",
                     18138 => "00101001",
                     18139 => "00000111",
                     18140 => "10101000",
                     18141 => "10111001",
                     18142 => "10010000",
                     18143 => "11000110",
                     18144 => "00101100",
                     18145 => "11011101",
                     18146 => "00000110",
                     18147 => "11110000",
                     18148 => "00000111",
                     18149 => "11001000",
                     18150 => "10011000",
                     18151 => "00101001",
                     18152 => "00000111",
                     18153 => "01001100",
                     18154 => "11011100",
                     18155 => "11000110",
                     18156 => "00001101",
                     18157 => "11011101",
                     18158 => "00000110",
                     18159 => "10001101",
                     18160 => "11011101",
                     18161 => "00000110",
                     18162 => "10111001",
                     18163 => "10011000",
                     18164 => "11000110",
                     18165 => "00100000",
                     18166 => "11011110",
                     18167 => "11000101",
                     18168 => "10011101",
                     18169 => "00010111",
                     18170 => "00000100",
                     18171 => "10101001",
                     18172 => "00100000",
                     18173 => "10001101",
                     18174 => "10001111",
                     18175 => "00000111",
                     18176 => "01001100",
                     18177 => "01110010",
                     18178 => "11000010",
                     18179 => "10100000",
                     18180 => "11111111",
                     18181 => "11001000",
                     18182 => "11000000",
                     18183 => "00000101",
                     18184 => "10110000",
                     18185 => "00001101",
                     18186 => "10111001",
                     18187 => "00001111",
                     18188 => "00000000",
                     18189 => "11110000",
                     18190 => "11110110",
                     18191 => "10111001",
                     18192 => "00010110",
                     18193 => "00000000",
                     18194 => "11001001",
                     18195 => "00001000",
                     18196 => "11010000",
                     18197 => "11101111",
                     18198 => "01100000",
                     18199 => "10100101",
                     18200 => "11111110",
                     18201 => "00001001",
                     18202 => "00001000",
                     18203 => "10000101",
                     18204 => "11111110",
                     18205 => "10101001",
                     18206 => "00001000",
                     18207 => "11010000",
                     18208 => "10101000",
                     18209 => "10100000",
                     18210 => "00000000",
                     18211 => "00111000",
                     18212 => "11101001",
                     18213 => "00110111",
                     18214 => "01001000",
                     18215 => "11001001",
                     18216 => "00000100",
                     18217 => "10110000",
                     18218 => "00001011",
                     18219 => "01001000",
                     18220 => "10100000",
                     18221 => "00000110",
                     18222 => "10101101",
                     18223 => "01101010",
                     18224 => "00000111",
                     18225 => "11110000",
                     18226 => "00000010",
                     18227 => "10100000",
                     18228 => "00000010",
                     18229 => "01101000",
                     18230 => "10000100",
                     18231 => "00000001",
                     18232 => "10100000",
                     18233 => "10110000",
                     18234 => "00101001",
                     18235 => "00000010",
                     18236 => "11110000",
                     18237 => "00000010",
                     18238 => "10100000",
                     18239 => "01110000",
                     18240 => "10000100",
                     18241 => "00000000",
                     18242 => "10101101",
                     18243 => "00011011",
                     18244 => "00000111",
                     18245 => "10000101",
                     18246 => "00000010",
                     18247 => "10101101",
                     18248 => "00011101",
                     18249 => "00000111",
                     18250 => "10000101",
                     18251 => "00000011",
                     18252 => "10100000",
                     18253 => "00000010",
                     18254 => "01101000",
                     18255 => "01001010",
                     18256 => "10010000",
                     18257 => "00000001",
                     18258 => "11001000",
                     18259 => "10001100",
                     18260 => "11010011",
                     18261 => "00000110",
                     18262 => "10100010",
                     18263 => "11111111",
                     18264 => "11101000",
                     18265 => "11100000",
                     18266 => "00000101",
                     18267 => "10110000",
                     18268 => "00101101",
                     18269 => "10110101",
                     18270 => "00001111",
                     18271 => "11010000",
                     18272 => "11110111",
                     18273 => "10100101",
                     18274 => "00000001",
                     18275 => "10010101",
                     18276 => "00010110",
                     18277 => "10100101",
                     18278 => "00000010",
                     18279 => "10010101",
                     18280 => "01101110",
                     18281 => "10100101",
                     18282 => "00000011",
                     18283 => "10010101",
                     18284 => "10000111",
                     18285 => "00011000",
                     18286 => "01101001",
                     18287 => "00011000",
                     18288 => "10000101",
                     18289 => "00000011",
                     18290 => "10100101",
                     18291 => "00000010",
                     18292 => "01101001",
                     18293 => "00000000",
                     18294 => "10000101",
                     18295 => "00000010",
                     18296 => "10100101",
                     18297 => "00000000",
                     18298 => "10010101",
                     18299 => "11001111",
                     18300 => "10101001",
                     18301 => "00000001",
                     18302 => "10010101",
                     18303 => "10110110",
                     18304 => "10010101",
                     18305 => "00001111",
                     18306 => "00100000",
                     18307 => "01110010",
                     18308 => "11000010",
                     18309 => "11001110",
                     18310 => "11010011",
                     18311 => "00000110",
                     18312 => "11010000",
                     18313 => "11001100",
                     18314 => "01001100",
                     18315 => "01100100",
                     18316 => "11000010",
                     18317 => "10101001",
                     18318 => "00000001",
                     18319 => "10010101",
                     18320 => "01011000",
                     18321 => "01001010",
                     18322 => "10010101",
                     18323 => "00011110",
                     18324 => "10010101",
                     18325 => "10100000",
                     18326 => "10110101",
                     18327 => "11001111",
                     18328 => "10011101",
                     18329 => "00110100",
                     18330 => "00000100",
                     18331 => "00111000",
                     18332 => "11101001",
                     18333 => "00011000",
                     18334 => "10011101",
                     18335 => "00010111",
                     18336 => "00000100",
                     18337 => "10101001",
                     18338 => "00001001",
                     18339 => "01001100",
                     18340 => "11100001",
                     18341 => "11000111",
                     18342 => "10110101",
                     18343 => "00010110",
                     18344 => "10001101",
                     18345 => "11001011",
                     18346 => "00000110",
                     18347 => "00111000",
                     18348 => "11101001",
                     18349 => "00010010",
                     18350 => "00100000",
                     18351 => "00000100",
                     18352 => "10001110",
                     18353 => "10101010",
                     18354 => "11000011",
                     18355 => "10111101",
                     18356 => "11000111",
                     18357 => "10101110",
                     18358 => "11000100",
                     18359 => "10101001",
                     18360 => "11000101",
                     18361 => "01000011",
                     18362 => "11000110",
                     18363 => "10100010",
                     18364 => "11000110",
                     18365 => "01100000",
                     18366 => "10100000",
                     18367 => "00000101",
                     18368 => "10111001",
                     18369 => "00010110",
                     18370 => "00000000",
                     18371 => "11001001",
                     18372 => "00010001",
                     18373 => "11010000",
                     18374 => "00000101",
                     18375 => "10101001",
                     18376 => "00000001",
                     18377 => "10011001",
                     18378 => "00011110",
                     18379 => "00000000",
                     18380 => "10001000",
                     18381 => "00010000",
                     18382 => "11110001",
                     18383 => "10101001",
                     18384 => "00000000",
                     18385 => "10001101",
                     18386 => "11001011",
                     18387 => "00000110",
                     18388 => "10010101",
                     18389 => "00001111",
                     18390 => "01100000",
                     18391 => "10101001",
                     18392 => "00000010",
                     18393 => "10010101",
                     18394 => "01000110",
                     18395 => "10101001",
                     18396 => "11110110",
                     18397 => "10010101",
                     18398 => "01011000",
                     18399 => "10101001",
                     18400 => "00000011",
                     18401 => "10011101",
                     18402 => "10011010",
                     18403 => "00000100",
                     18404 => "01100000",
                     18405 => "11010110",
                     18406 => "11001111",
                     18407 => "11010110",
                     18408 => "11001111",
                     18409 => "10101100",
                     18410 => "11001100",
                     18411 => "00000110",
                     18412 => "11010000",
                     18413 => "00000101",
                     18414 => "10100000",
                     18415 => "00000010",
                     18416 => "00100000",
                     18417 => "01110111",
                     18418 => "11001000",
                     18419 => "10100000",
                     18420 => "11111111",
                     18421 => "10101101",
                     18422 => "10100000",
                     18423 => "00000011",
                     18424 => "10010101",
                     18425 => "00011110",
                     18426 => "00010000",
                     18427 => "00000010",
                     18428 => "10001010",
                     18429 => "10101000",
                     18430 => "10001100",
                     18431 => "10100000",
                     18432 => "00000011",
                     18433 => "10101001",
                     18434 => "00000000",
                     18435 => "10010101",
                     18436 => "01000110",
                     18437 => "10101000",
                     18438 => "00100000",
                     18439 => "01110111",
                     18440 => "11001000",
                     18441 => "10101001",
                     18442 => "11111111",
                     18443 => "10011101",
                     18444 => "10100010",
                     18445 => "00000011",
                     18446 => "01001100",
                     18447 => "00101110",
                     18448 => "11001000",
                     18449 => "10101001",
                     18450 => "00000000",
                     18451 => "10010101",
                     18452 => "01011000",
                     18453 => "01001100",
                     18454 => "00101110",
                     18455 => "11001000",
                     18456 => "10100000",
                     18457 => "01000000",
                     18458 => "10110101",
                     18459 => "11001111",
                     18460 => "00010000",
                     18461 => "00000111",
                     18462 => "01001001",
                     18463 => "11111111",
                     18464 => "00011000",
                     18465 => "01101001",
                     18466 => "00000001",
                     18467 => "10100000",
                     18468 => "11000000",
                     18469 => "10011101",
                     18470 => "00000001",
                     18471 => "00000100",
                     18472 => "10011000",
                     18473 => "00011000",
                     18474 => "01110101",
                     18475 => "11001111",
                     18476 => "10010101",
                     18477 => "01011000",
                     18478 => "00100000",
                     18479 => "01101001",
                     18480 => "11000011",
                     18481 => "10101001",
                     18482 => "00000101",
                     18483 => "10101100",
                     18484 => "01001110",
                     18485 => "00000111",
                     18486 => "11000000",
                     18487 => "00000011",
                     18488 => "11110000",
                     18489 => "00000111",
                     18490 => "10101100",
                     18491 => "11001100",
                     18492 => "00000110",
                     18493 => "11010000",
                     18494 => "00000010",
                     18495 => "10101001",
                     18496 => "00000110",
                     18497 => "10011101",
                     18498 => "10011010",
                     18499 => "00000100",
                     18500 => "01100000",
                     18501 => "00100000",
                     18502 => "01010001",
                     18503 => "11001000",
                     18504 => "01001100",
                     18505 => "01001110",
                     18506 => "11001000",
                     18507 => "00100000",
                     18508 => "01011101",
                     18509 => "11001000",
                     18510 => "01001100",
                     18511 => "00110001",
                     18512 => "11001000",
                     18513 => "10101001",
                     18514 => "00010000",
                     18515 => "10011101",
                     18516 => "00110100",
                     18517 => "00000100",
                     18518 => "10101001",
                     18519 => "11111111",
                     18520 => "10010101",
                     18521 => "10100000",
                     18522 => "01001100",
                     18523 => "01100110",
                     18524 => "11001000",
                     18525 => "10101001",
                     18526 => "11110000",
                     18527 => "10011101",
                     18528 => "00110100",
                     18529 => "00000100",
                     18530 => "10101001",
                     18531 => "00000000",
                     18532 => "10010101",
                     18533 => "10100000",
                     18534 => "10100000",
                     18535 => "00000001",
                     18536 => "00100000",
                     18537 => "01110111",
                     18538 => "11001000",
                     18539 => "10101001",
                     18540 => "00000100",
                     18541 => "10011101",
                     18542 => "10011010",
                     18543 => "00000100",
                     18544 => "01100000",
                     18545 => "00001000",
                     18546 => "00001100",
                     18547 => "11111000",
                     18548 => "00000000",
                     18549 => "00000000",
                     18550 => "11111111",
                     18551 => "10110101",
                     18552 => "10000111",
                     18553 => "00011000",
                     18554 => "01111001",
                     18555 => "01110001",
                     18556 => "11001000",
                     18557 => "10010101",
                     18558 => "10000111",
                     18559 => "10110101",
                     18560 => "01101110",
                     18561 => "01111001",
                     18562 => "01110100",
                     18563 => "11001000",
                     18564 => "10010101",
                     18565 => "01101110",
                     18566 => "01100000",
                     18567 => "01100000",
                     18568 => "10100110",
                     18569 => "00001000",
                     18570 => "10101001",
                     18571 => "00000000",
                     18572 => "10110100",
                     18573 => "00010110",
                     18574 => "11000000",
                     18575 => "00010101",
                     18576 => "10010000",
                     18577 => "00000011",
                     18578 => "10011000",
                     18579 => "11101001",
                     18580 => "00010100",
                     18581 => "00100000",
                     18582 => "00000100",
                     18583 => "10001110",
                     18584 => "11100110",
                     18585 => "11001000",
                     18586 => "00111011",
                     18587 => "11001001",
                     18588 => "01011101",
                     18589 => "11010010",
                     18590 => "11011100",
                     18591 => "11001000",
                     18592 => "11011100",
                     18593 => "11001000",
                     18594 => "11011100",
                     18595 => "11001000",
                     18596 => "11011100",
                     18597 => "11001000",
                     18598 => "01001101",
                     18599 => "11001001",
                     18600 => "01001101",
                     18601 => "11001001",
                     18602 => "01001101",
                     18603 => "11001001",
                     18604 => "01001101",
                     18605 => "11001001",
                     18606 => "01001101",
                     18607 => "11001001",
                     18608 => "01001101",
                     18609 => "11001001",
                     18610 => "01001101",
                     18611 => "11001001",
                     18612 => "01001101",
                     18613 => "11001001",
                     18614 => "11011100",
                     18615 => "11001000",
                     18616 => "01101011",
                     18617 => "11001001",
                     18618 => "01101011",
                     18619 => "11001001",
                     18620 => "01101011",
                     18621 => "11001001",
                     18622 => "01101011",
                     18623 => "11001001",
                     18624 => "01101011",
                     18625 => "11001001",
                     18626 => "01101011",
                     18627 => "11001001",
                     18628 => "01101011",
                     18629 => "11001001",
                     18630 => "01010011",
                     18631 => "11001001",
                     18632 => "01010011",
                     18633 => "11001001",
                     18634 => "00101101",
                     18635 => "11010000",
                     18636 => "10001010",
                     18637 => "10111100",
                     18638 => "01010000",
                     18639 => "10111001",
                     18640 => "11011100",
                     18641 => "11001000",
                     18642 => "10100001",
                     18643 => "11010010",
                     18644 => "10111010",
                     18645 => "10111000",
                     18646 => "11011100",
                     18647 => "11001000",
                     18648 => "10100100",
                     18649 => "10110111",
                     18650 => "11011101",
                     18651 => "11001000",
                     18652 => "01100000",
                     18653 => "00100000",
                     18654 => "10110110",
                     18655 => "11110001",
                     18656 => "00100000",
                     18657 => "01011001",
                     18658 => "11110001",
                     18659 => "01001100",
                     18660 => "10000100",
                     18661 => "11101000",
                     18662 => "10101001",
                     18663 => "00000000",
                     18664 => "10011101",
                     18665 => "11000101",
                     18666 => "00000011",
                     18667 => "00100000",
                     18668 => "10110110",
                     18669 => "11110001",
                     18670 => "00100000",
                     18671 => "01011001",
                     18672 => "11110001",
                     18673 => "00100000",
                     18674 => "10000100",
                     18675 => "11101000",
                     18676 => "00100000",
                     18677 => "01001011",
                     18678 => "11100010",
                     18679 => "00100000",
                     18680 => "11001001",
                     18681 => "11011111",
                     18682 => "00100000",
                     18683 => "00110101",
                     18684 => "11011010",
                     18685 => "00100000",
                     18686 => "01010011",
                     18687 => "11011000",
                     18688 => "10101100",
                     18689 => "01000111",
                     18690 => "00000111",
                     18691 => "11010000",
                     18692 => "00000011",
                     18693 => "00100000",
                     18694 => "00001011",
                     18695 => "11001001",
                     18696 => "01001100",
                     18697 => "01000010",
                     18698 => "11010110",
                     18699 => "10110101",
                     18700 => "00010110",
                     18701 => "00100000",
                     18702 => "00000100",
                     18703 => "10001110",
                     18704 => "01111101",
                     18705 => "11001010",
                     18706 => "01111101",
                     18707 => "11001010",
                     18708 => "01111101",
                     18709 => "11001010",
                     18710 => "01111101",
                     18711 => "11001010",
                     18712 => "01111101",
                     18713 => "11001010",
                     18714 => "11011110",
                     18715 => "11001001",
                     18716 => "01111101",
                     18717 => "11001010",
                     18718 => "10001111",
                     18719 => "11001011",
                     18720 => "00111100",
                     18721 => "11001100",
                     18722 => "00111010",
                     18723 => "11001001",
                     18724 => "01010000",
                     18725 => "11001100",
                     18726 => "01010000",
                     18727 => "11001100",
                     18728 => "10110110",
                     18729 => "11001001",
                     18730 => "01111000",
                     18731 => "11010011",
                     18732 => "11111111",
                     18733 => "11001010",
                     18734 => "00000101",
                     18735 => "11001011",
                     18736 => "00101011",
                     18737 => "11001011",
                     18738 => "11110000",
                     18739 => "11001110",
                     18740 => "01111101",
                     18741 => "11001010",
                     18742 => "00111010",
                     18743 => "11001001",
                     18744 => "11011011",
                     18745 => "11001110",
                     18746 => "01100000",
                     18747 => "00100000",
                     18748 => "10110011",
                     18749 => "11010001",
                     18750 => "00100000",
                     18751 => "10110110",
                     18752 => "11110001",
                     18753 => "00100000",
                     18754 => "01011001",
                     18755 => "11110001",
                     18756 => "00100000",
                     18757 => "01001011",
                     18758 => "11100010",
                     18759 => "00100000",
                     18760 => "01010011",
                     18761 => "11011000",
                     18762 => "01001100",
                     18763 => "01000010",
                     18764 => "11010110",
                     18765 => "00100000",
                     18766 => "01000010",
                     18767 => "11001101",
                     18768 => "01001100",
                     18769 => "01000010",
                     18770 => "11010110",
                     18771 => "00100000",
                     18772 => "10110110",
                     18773 => "11110001",
                     18774 => "00100000",
                     18775 => "01011001",
                     18776 => "11110001",
                     18777 => "00100000",
                     18778 => "01010100",
                     18779 => "11100010",
                     18780 => "00100000",
                     18781 => "01111101",
                     18782 => "11011011",
                     18783 => "00100000",
                     18784 => "01011001",
                     18785 => "11110001",
                     18786 => "00100000",
                     18787 => "01101101",
                     18788 => "11101101",
                     18789 => "00100000",
                     18790 => "00011101",
                     18791 => "11010110",
                     18792 => "01001100",
                     18793 => "01000010",
                     18794 => "11010110",
                     18795 => "00100000",
                     18796 => "10110110",
                     18797 => "11110001",
                     18798 => "00100000",
                     18799 => "01011001",
                     18800 => "11110001",
                     18801 => "00100000",
                     18802 => "01111011",
                     18803 => "11100010",
                     18804 => "00100000",
                     18805 => "01000111",
                     18806 => "11011011",
                     18807 => "10101101",
                     18808 => "01000111",
                     18809 => "00000111",
                     18810 => "11010000",
                     18811 => "00000011",
                     18812 => "00100000",
                     18813 => "10001000",
                     18814 => "11001001",
                     18815 => "00100000",
                     18816 => "01011001",
                     18817 => "11110001",
                     18818 => "00100000",
                     18819 => "11001111",
                     18820 => "11100101",
                     18821 => "01001100",
                     18822 => "01000010",
                     18823 => "11010110",
                     18824 => "10110101",
                     18825 => "00010110",
                     18826 => "00111000",
                     18827 => "11101001",
                     18828 => "00100100",
                     18829 => "00100000",
                     18830 => "00000100",
                     18831 => "10001110",
                     18832 => "11111010",
                     18833 => "11010011",
                     18834 => "10011011",
                     18835 => "11010101",
                     18836 => "00010111",
                     18837 => "11010110",
                     18838 => "00010111",
                     18839 => "11010110",
                     18840 => "11001111",
                     18841 => "11010101",
                     18842 => "11111001",
                     18843 => "11010101",
                     18844 => "00000101",
                     18845 => "11010110",
                     18846 => "10101001",
                     18847 => "00000000",
                     18848 => "10010101",
                     18849 => "00001111",
                     18850 => "10010101",
                     18851 => "00010110",
                     18852 => "10010101",
                     18853 => "00011110",
                     18854 => "10011101",
                     18855 => "00010000",
                     18856 => "00000001",
                     18857 => "10011101",
                     18858 => "10010110",
                     18859 => "00000111",
                     18860 => "10011101",
                     18861 => "00100101",
                     18862 => "00000001",
                     18863 => "10011101",
                     18864 => "11000101",
                     18865 => "00000011",
                     18866 => "10011101",
                     18867 => "10001010",
                     18868 => "00000111",
                     18869 => "01100000",
                     18870 => "10111101",
                     18871 => "10010110",
                     18872 => "00000111",
                     18873 => "11010000",
                     18874 => "00010110",
                     18875 => "00100000",
                     18876 => "11111101",
                     18877 => "11000010",
                     18878 => "10111101",
                     18879 => "10101000",
                     18880 => "00000111",
                     18881 => "00001001",
                     18882 => "10000000",
                     18883 => "10011101",
                     18884 => "00110100",
                     18885 => "00000100",
                     18886 => "00101001",
                     18887 => "00001111",
                     18888 => "00001001",
                     18889 => "00000110",
                     18890 => "10011101",
                     18891 => "10010110",
                     18892 => "00000111",
                     18893 => "10101001",
                     18894 => "11111001",
                     18895 => "10010101",
                     18896 => "10100000",
                     18897 => "01001100",
                     18898 => "10010111",
                     18899 => "10111111",
                     18900 => "00110000",
                     18901 => "00011100",
                     18902 => "00000000",
                     18903 => "11101000",
                     18904 => "00000000",
                     18905 => "00011000",
                     18906 => "00001000",
                     18907 => "11111000",
                     18908 => "00001100",
                     18909 => "11110100",
                     18910 => "10110101",
                     18911 => "00011110",
                     18912 => "00101001",
                     18913 => "00100000",
                     18914 => "11110000",
                     18915 => "00000011",
                     18916 => "01001100",
                     18917 => "11101011",
                     18918 => "11001010",
                     18919 => "10110101",
                     18920 => "00111100",
                     18921 => "11110000",
                     18922 => "00101101",
                     18923 => "11010110",
                     18924 => "00111100",
                     18925 => "10101101",
                     18926 => "11010001",
                     18927 => "00000011",
                     18928 => "00101001",
                     18929 => "00001100",
                     18930 => "11010000",
                     18931 => "01101010",
                     18932 => "10111101",
                     18933 => "10100010",
                     18934 => "00000011",
                     18935 => "11010000",
                     18936 => "00010111",
                     18937 => "10101100",
                     18938 => "11001100",
                     18939 => "00000110",
                     18940 => "10111001",
                     18941 => "11010100",
                     18942 => "11001001",
                     18943 => "10011101",
                     18944 => "10100010",
                     18945 => "00000011",
                     18946 => "00100000",
                     18947 => "10011001",
                     18948 => "10111010",
                     18949 => "10010000",
                     18950 => "00001001",
                     18951 => "10110101",
                     18952 => "00011110",
                     18953 => "00001001",
                     18954 => "00001000",
                     18955 => "10010101",
                     18956 => "00011110",
                     18957 => "01001100",
                     18958 => "01011110",
                     18959 => "11001010",
                     18960 => "11011110",
                     18961 => "10100010",
                     18962 => "00000011",
                     18963 => "01001100",
                     18964 => "01011110",
                     18965 => "11001010",
                     18966 => "00100000",
                     18967 => "00110111",
                     18968 => "10110101",
                     18969 => "00011110",
                     18970 => "00101001",
                     18971 => "00000111",
                     18972 => "11001001",
                     18973 => "00000001",
                     18974 => "11110000",
                     18975 => "00111110",
                     18976 => "10101001",
                     18977 => "00000000",
                     18978 => "10000101",
                     18979 => "00000000",
                     18980 => "10100000",
                     18981 => "11111010",
                     18982 => "10110101",
                     18983 => "11001111",
                     18984 => "00110000",
                     18985 => "00010011",
                     18986 => "10100000",
                     18987 => "11111101",
                     18988 => "11001001",
                     18989 => "01110000",
                     18990 => "11100110",
                     18991 => "00000000",
                     18992 => "10010000",
                     18993 => "00001011",
                     18994 => "11000110",
                     18995 => "00000000",
                     18996 => "10111101",
                     18997 => "10101000",
                     18998 => "00000111",
                     18999 => "00101001",
                     19000 => "00000001",
                     19001 => "11010000",
                     19002 => "00000010",
                     19003 => "10100000",
                     19004 => "11111010",
                     19005 => "10010100",
                     19006 => "10100000",
                     19007 => "10110101",
                     19008 => "00011110",
                     19009 => "00001001",
                     19010 => "00000001",
                     19011 => "10010101",
                     19012 => "00011110",
                     19013 => "10100101",
                     19014 => "00000000",
                     19015 => "00111101",
                     19016 => "10101001",
                     19017 => "00000111",
                     19018 => "10101000",
                     19019 => "10101101",
                     19020 => "11001100",
                     19021 => "00000110",
                     19022 => "11010000",
                     19023 => "00000001",
                     19024 => "10101000",
                     19025 => "10111001",
                     19026 => "00010110",
                     19027 => "11001010",
                     19028 => "10011101",
                     19029 => "10001010",
                     19030 => "00000111",
                     19031 => "10111101",
                     19032 => "10101000",
                     19033 => "00000111",
                     19034 => "00001001",
                     19035 => "11000000",
                     19036 => "10010101",
                     19037 => "00111100",
                     19038 => "10100000",
                     19039 => "11111011",
                     19040 => "10100101",
                     19041 => "00001001",
                     19042 => "00101001",
                     19043 => "01000000",
                     19044 => "11010000",
                     19045 => "00000010",
                     19046 => "10100000",
                     19047 => "00000101",
                     19048 => "10010100",
                     19049 => "01011000",
                     19050 => "10100000",
                     19051 => "00000001",
                     19052 => "00100000",
                     19053 => "01001011",
                     19054 => "11100001",
                     19055 => "00110000",
                     19056 => "00001010",
                     19057 => "11001000",
                     19058 => "10111101",
                     19059 => "10010110",
                     19060 => "00000111",
                     19061 => "11010000",
                     19062 => "00000100",
                     19063 => "10101001",
                     19064 => "11110110",
                     19065 => "10010101",
                     19066 => "01011000",
                     19067 => "10010100",
                     19068 => "01000110",
                     19069 => "10100000",
                     19070 => "00000000",
                     19071 => "10110101",
                     19072 => "00011110",
                     19073 => "00101001",
                     19074 => "01000000",
                     19075 => "11010000",
                     19076 => "00011001",
                     19077 => "10110101",
                     19078 => "00011110",
                     19079 => "00001010",
                     19080 => "10110000",
                     19081 => "00110000",
                     19082 => "10110101",
                     19083 => "00011110",
                     19084 => "00101001",
                     19085 => "00100000",
                     19086 => "11010000",
                     19087 => "01011011",
                     19088 => "10110101",
                     19089 => "00011110",
                     19090 => "00101001",
                     19091 => "00000111",
                     19092 => "11110000",
                     19093 => "00100100",
                     19094 => "11001001",
                     19095 => "00000101",
                     19096 => "11110000",
                     19097 => "00000100",
                     19098 => "11001001",
                     19099 => "00000011",
                     19100 => "10110000",
                     19101 => "00110000",
                     19102 => "00100000",
                     19103 => "01101000",
                     19104 => "10111111",
                     19105 => "10100000",
                     19106 => "00000000",
                     19107 => "10110101",
                     19108 => "00011110",
                     19109 => "11001001",
                     19110 => "00000010",
                     19111 => "11110000",
                     19112 => "00001100",
                     19113 => "00101001",
                     19114 => "01000000",
                     19115 => "11110000",
                     19116 => "00001101",
                     19117 => "10110101",
                     19118 => "00010110",
                     19119 => "11001001",
                     19120 => "00101110",
                     19121 => "11110000",
                     19122 => "00000111",
                     19123 => "11010000",
                     19124 => "00000011",
                     19125 => "01001100",
                     19126 => "00000111",
                     19127 => "10111111",
                     19128 => "10100000",
                     19129 => "00000001",
                     19130 => "10110101",
                     19131 => "01011000",
                     19132 => "01001000",
                     19133 => "00010000",
                     19134 => "00000010",
                     19135 => "11001000",
                     19136 => "11001000",
                     19137 => "00011000",
                     19138 => "01111001",
                     19139 => "11010110",
                     19140 => "11001001",
                     19141 => "10010101",
                     19142 => "01011000",
                     19143 => "00100000",
                     19144 => "00000111",
                     19145 => "10111111",
                     19146 => "01101000",
                     19147 => "10010101",
                     19148 => "01011000",
                     19149 => "01100000",
                     19150 => "10111101",
                     19151 => "10010110",
                     19152 => "00000111",
                     19153 => "11010000",
                     19154 => "00011110",
                     19155 => "10010101",
                     19156 => "00011110",
                     19157 => "10100101",
                     19158 => "00001001",
                     19159 => "00101001",
                     19160 => "00000001",
                     19161 => "10101000",
                     19162 => "11001000",
                     19163 => "10010100",
                     19164 => "01000110",
                     19165 => "10001000",
                     19166 => "10101101",
                     19167 => "01101010",
                     19168 => "00000111",
                     19169 => "11110000",
                     19170 => "00000010",
                     19171 => "11001000",
                     19172 => "11001000",
                     19173 => "10111001",
                     19174 => "11011010",
                     19175 => "11001001",
                     19176 => "10010101",
                     19177 => "01011000",
                     19178 => "01100000",
                     19179 => "00100000",
                     19180 => "01101000",
                     19181 => "10111111",
                     19182 => "01001100",
                     19183 => "00000111",
                     19184 => "10111111",
                     19185 => "11001001",
                     19186 => "00001011",
                     19187 => "11010000",
                     19188 => "00001001",
                     19189 => "10110101",
                     19190 => "00010110",
                     19191 => "11001001",
                     19192 => "00000110",
                     19193 => "11010000",
                     19194 => "00000011",
                     19195 => "00100000",
                     19196 => "10011110",
                     19197 => "11001001",
                     19198 => "01100000",
                     19199 => "00100000",
                     19200 => "10010111",
                     19201 => "10111111",
                     19202 => "01001100",
                     19203 => "00000111",
                     19204 => "10111111",
                     19205 => "10110101",
                     19206 => "10100000",
                     19207 => "00011101",
                     19208 => "00110100",
                     19209 => "00000100",
                     19210 => "11010000",
                     19211 => "00010011",
                     19212 => "10011101",
                     19213 => "00010111",
                     19214 => "00000100",
                     19215 => "10110101",
                     19216 => "11001111",
                     19217 => "11011101",
                     19218 => "00000001",
                     19219 => "00000100",
                     19220 => "10110000",
                     19221 => "00001001",
                     19222 => "10100101",
                     19223 => "00001001",
                     19224 => "00101001",
                     19225 => "00000111",
                     19226 => "11010000",
                     19227 => "00000010",
                     19228 => "11110110",
                     19229 => "11001111",
                     19230 => "01100000",
                     19231 => "10110101",
                     19232 => "11001111",
                     19233 => "11010101",
                     19234 => "01011000",
                     19235 => "10010000",
                     19236 => "00000011",
                     19237 => "01001100",
                     19238 => "01111010",
                     19239 => "10111111",
                     19240 => "01001100",
                     19241 => "01110101",
                     19242 => "10111111",
                     19243 => "00100000",
                     19244 => "01001011",
                     19245 => "11001011",
                     19246 => "00100000",
                     19247 => "01101100",
                     19248 => "11001011",
                     19249 => "10100000",
                     19250 => "00000001",
                     19251 => "10100101",
                     19252 => "00001001",
                     19253 => "00101001",
                     19254 => "00000011",
                     19255 => "11010000",
                     19256 => "00010001",
                     19257 => "10100101",
                     19258 => "00001001",
                     19259 => "00101001",
                     19260 => "01000000",
                     19261 => "11010000",
                     19262 => "00000010",
                     19263 => "10100000",
                     19264 => "11111111",
                     19265 => "10000100",
                     19266 => "00000000",
                     19267 => "10110101",
                     19268 => "11001111",
                     19269 => "00011000",
                     19270 => "01100101",
                     19271 => "00000000",
                     19272 => "10010101",
                     19273 => "11001111",
                     19274 => "01100000",
                     19275 => "10101001",
                     19276 => "00010011",
                     19277 => "10000101",
                     19278 => "00000001",
                     19279 => "10100101",
                     19280 => "00001001",
                     19281 => "00101001",
                     19282 => "00000011",
                     19283 => "11010000",
                     19284 => "00001101",
                     19285 => "10110100",
                     19286 => "01011000",
                     19287 => "10110101",
                     19288 => "10100000",
                     19289 => "01001010",
                     19290 => "10110000",
                     19291 => "00001010",
                     19292 => "11000100",
                     19293 => "00000001",
                     19294 => "11110000",
                     19295 => "00000011",
                     19296 => "11110110",
                     19297 => "01011000",
                     19298 => "01100000",
                     19299 => "11110110",
                     19300 => "10100000",
                     19301 => "01100000",
                     19302 => "10011000",
                     19303 => "11110000",
                     19304 => "11111010",
                     19305 => "11010110",
                     19306 => "01011000",
                     19307 => "01100000",
                     19308 => "10110101",
                     19309 => "01011000",
                     19310 => "01001000",
                     19311 => "10100000",
                     19312 => "00000001",
                     19313 => "10110101",
                     19314 => "10100000",
                     19315 => "00101001",
                     19316 => "00000010",
                     19317 => "11010000",
                     19318 => "00001011",
                     19319 => "10110101",
                     19320 => "01011000",
                     19321 => "01001001",
                     19322 => "11111111",
                     19323 => "00011000",
                     19324 => "01101001",
                     19325 => "00000001",
                     19326 => "10010101",
                     19327 => "01011000",
                     19328 => "10100000",
                     19329 => "00000010",
                     19330 => "10010100",
                     19331 => "01000110",
                     19332 => "00100000",
                     19333 => "00000111",
                     19334 => "10111111",
                     19335 => "10000101",
                     19336 => "00000000",
                     19337 => "01101000",
                     19338 => "10010101",
                     19339 => "01011000",
                     19340 => "01100000",
                     19341 => "00000111",
                     19342 => "00000001",
                     19343 => "10110101",
                     19344 => "00011110",
                     19345 => "00101001",
                     19346 => "00100000",
                     19347 => "11010000",
                     19348 => "01001101",
                     19349 => "10101100",
                     19350 => "11001100",
                     19351 => "00000110",
                     19352 => "10111101",
                     19353 => "10101000",
                     19354 => "00000111",
                     19355 => "00111001",
                     19356 => "10001101",
                     19357 => "11001011",
                     19358 => "11010000",
                     19359 => "00010010",
                     19360 => "10001010",
                     19361 => "01001010",
                     19362 => "10010000",
                     19363 => "00000100",
                     19364 => "10100100",
                     19365 => "01000101",
                     19366 => "10110000",
                     19367 => "00001000",
                     19368 => "10100000",
                     19369 => "00000010",
                     19370 => "00100000",
                     19371 => "01001011",
                     19372 => "11100001",
                     19373 => "00010000",
                     19374 => "00000001",
                     19375 => "10001000",
                     19376 => "10010100",
                     19377 => "01000110",
                     19378 => "00100000",
                     19379 => "11100101",
                     19380 => "11001011",
                     19381 => "10110101",
                     19382 => "11001111",
                     19383 => "00111000",
                     19384 => "11111101",
                     19385 => "00110100",
                     19386 => "00000100",
                     19387 => "11001001",
                     19388 => "00100000",
                     19389 => "10010000",
                     19390 => "00000010",
                     19391 => "10010101",
                     19392 => "11001111",
                     19393 => "10110100",
                     19394 => "01000110",
                     19395 => "10001000",
                     19396 => "11010000",
                     19397 => "00001110",
                     19398 => "10110101",
                     19399 => "10000111",
                     19400 => "00011000",
                     19401 => "01110101",
                     19402 => "01011000",
                     19403 => "10010101",
                     19404 => "10000111",
                     19405 => "10110101",
                     19406 => "01101110",
                     19407 => "01101001",
                     19408 => "00000000",
                     19409 => "10010101",
                     19410 => "01101110",
                     19411 => "01100000",
                     19412 => "10110101",
                     19413 => "10000111",
                     19414 => "00111000",
                     19415 => "11110101",
                     19416 => "01011000",
                     19417 => "10010101",
                     19418 => "10000111",
                     19419 => "10110101",
                     19420 => "01101110",
                     19421 => "11101001",
                     19422 => "00000000",
                     19423 => "10010101",
                     19424 => "01101110",
                     19425 => "01100000",
                     19426 => "01001100",
                     19427 => "10010001",
                     19428 => "10111111",
                     19429 => "10110101",
                     19430 => "10100000",
                     19431 => "00101001",
                     19432 => "00000010",
                     19433 => "11010000",
                     19434 => "00110111",
                     19435 => "10100101",
                     19436 => "00001001",
                     19437 => "00101001",
                     19438 => "00000111",
                     19439 => "01001000",
                     19440 => "10110101",
                     19441 => "10100000",
                     19442 => "01001010",
                     19443 => "10110000",
                     19444 => "00010101",
                     19445 => "01101000",
                     19446 => "11010000",
                     19447 => "00010001",
                     19448 => "10111101",
                     19449 => "00110100",
                     19450 => "00000100",
                     19451 => "00011000",
                     19452 => "01101001",
                     19453 => "00000001",
                     19454 => "10011101",
                     19455 => "00110100",
                     19456 => "00000100",
                     19457 => "10010101",
                     19458 => "01011000",
                     19459 => "11001001",
                     19460 => "00000010",
                     19461 => "11010000",
                     19462 => "00000010",
                     19463 => "11110110",
                     19464 => "10100000",
                     19465 => "01100000",
                     19466 => "01101000",
                     19467 => "11010000",
                     19468 => "00010100",
                     19469 => "10111101",
                     19470 => "00110100",
                     19471 => "00000100",
                     19472 => "00111000",
                     19473 => "11101001",
                     19474 => "00000001",
                     19475 => "10011101",
                     19476 => "00110100",
                     19477 => "00000100",
                     19478 => "10010101",
                     19479 => "01011000",
                     19480 => "11010000",
                     19481 => "00000111",
                     19482 => "11110110",
                     19483 => "10100000",
                     19484 => "10101001",
                     19485 => "00000010",
                     19486 => "10011101",
                     19487 => "10010110",
                     19488 => "00000111",
                     19489 => "01100000",
                     19490 => "10111101",
                     19491 => "10010110",
                     19492 => "00000111",
                     19493 => "11110000",
                     19494 => "00001000",
                     19495 => "10100101",
                     19496 => "00001001",
                     19497 => "01001010",
                     19498 => "10110000",
                     19499 => "00000010",
                     19500 => "11110110",
                     19501 => "11001111",
                     19502 => "01100000",
                     19503 => "10110101",
                     19504 => "11001111",
                     19505 => "01101001",
                     19506 => "00001100",
                     19507 => "11000101",
                     19508 => "11001110",
                     19509 => "10010000",
                     19510 => "11110000",
                     19511 => "10101001",
                     19512 => "00000000",
                     19513 => "10010101",
                     19514 => "10100000",
                     19515 => "01100000",
                     19516 => "10110101",
                     19517 => "00011110",
                     19518 => "00101001",
                     19519 => "00100000",
                     19520 => "11110000",
                     19521 => "00000011",
                     19522 => "01001100",
                     19523 => "10010111",
                     19524 => "10111111",
                     19525 => "10101001",
                     19526 => "11101000",
                     19527 => "10010101",
                     19528 => "01011000",
                     19529 => "01001100",
                     19530 => "00000111",
                     19531 => "10111111",
                     19532 => "01000000",
                     19533 => "10000000",
                     19534 => "00000100",
                     19535 => "00000100",
                     19536 => "10110101",
                     19537 => "00011110",
                     19538 => "00101001",
                     19539 => "00100000",
                     19540 => "11110000",
                     19541 => "00000011",
                     19542 => "01001100",
                     19543 => "10010001",
                     19544 => "10111111",
                     19545 => "10000101",
                     19546 => "00000011",
                     19547 => "10110101",
                     19548 => "00010110",
                     19549 => "00111000",
                     19550 => "11101001",
                     19551 => "00001010",
                     19552 => "10101000",
                     19553 => "10111001",
                     19554 => "01001100",
                     19555 => "11001100",
                     19556 => "10000101",
                     19557 => "00000010",
                     19558 => "10111101",
                     19559 => "00000001",
                     19560 => "00000100",
                     19561 => "00111000",
                     19562 => "11100101",
                     19563 => "00000010",
                     19564 => "10011101",
                     19565 => "00000001",
                     19566 => "00000100",
                     19567 => "10110101",
                     19568 => "10000111",
                     19569 => "11101001",
                     19570 => "00000000",
                     19571 => "10010101",
                     19572 => "10000111",
                     19573 => "10110101",
                     19574 => "01101110",
                     19575 => "11101001",
                     19576 => "00000000",
                     19577 => "10010101",
                     19578 => "01101110",
                     19579 => "10101001",
                     19580 => "00100000",
                     19581 => "10000101",
                     19582 => "00000010",
                     19583 => "11100000",
                     19584 => "00000010",
                     19585 => "10010000",
                     19586 => "01001001",
                     19587 => "10110101",
                     19588 => "01011000",
                     19589 => "11001001",
                     19590 => "00010000",
                     19591 => "10010000",
                     19592 => "00010110",
                     19593 => "10111101",
                     19594 => "00010111",
                     19595 => "00000100",
                     19596 => "00011000",
                     19597 => "01100101",
                     19598 => "00000010",
                     19599 => "10011101",
                     19600 => "00010111",
                     19601 => "00000100",
                     19602 => "10110101",
                     19603 => "11001111",
                     19604 => "01100101",
                     19605 => "00000011",
                     19606 => "10010101",
                     19607 => "11001111",
                     19608 => "10110101",
                     19609 => "10110110",
                     19610 => "01101001",
                     19611 => "00000000",
                     19612 => "01001100",
                     19613 => "10110010",
                     19614 => "11001100",
                     19615 => "10111101",
                     19616 => "00010111",
                     19617 => "00000100",
                     19618 => "00111000",
                     19619 => "11100101",
                     19620 => "00000010",
                     19621 => "10011101",
                     19622 => "00010111",
                     19623 => "00000100",
                     19624 => "10110101",
                     19625 => "11001111",
                     19626 => "11100101",
                     19627 => "00000011",
                     19628 => "10010101",
                     19629 => "11001111",
                     19630 => "10110101",
                     19631 => "10110110",
                     19632 => "11101001",
                     19633 => "00000000",
                     19634 => "10010101",
                     19635 => "10110110",
                     19636 => "10100000",
                     19637 => "00000000",
                     19638 => "10110101",
                     19639 => "11001111",
                     19640 => "00111000",
                     19641 => "11111101",
                     19642 => "00110100",
                     19643 => "00000100",
                     19644 => "00010000",
                     19645 => "00000111",
                     19646 => "10100000",
                     19647 => "00010000",
                     19648 => "01001001",
                     19649 => "11111111",
                     19650 => "00011000",
                     19651 => "01101001",
                     19652 => "00000001",
                     19653 => "11001001",
                     19654 => "00001111",
                     19655 => "10010000",
                     19656 => "00000011",
                     19657 => "10011000",
                     19658 => "10010101",
                     19659 => "01011000",
                     19660 => "01100000",
                     19661 => "00000000",
                     19662 => "00000001",
                     19663 => "00000011",
                     19664 => "00000100",
                     19665 => "00000101",
                     19666 => "00000110",
                     19667 => "00000111",
                     19668 => "00000111",
                     19669 => "00001000",
                     19670 => "00000000",
                     19671 => "00000011",
                     19672 => "00000110",
                     19673 => "00001001",
                     19674 => "00001011",
                     19675 => "00001101",
                     19676 => "00001110",
                     19677 => "00001111",
                     19678 => "00010000",
                     19679 => "00000000",
                     19680 => "00000100",
                     19681 => "00001001",
                     19682 => "00001101",
                     19683 => "00010000",
                     19684 => "00010011",
                     19685 => "00010110",
                     19686 => "00010111",
                     19687 => "00011000",
                     19688 => "00000000",
                     19689 => "00000110",
                     19690 => "00001100",
                     19691 => "00010010",
                     19692 => "00010110",
                     19693 => "00011010",
                     19694 => "00011101",
                     19695 => "00011111",
                     19696 => "00100000",
                     19697 => "00000000",
                     19698 => "00000111",
                     19699 => "00001111",
                     19700 => "00010110",
                     19701 => "00011100",
                     19702 => "00100001",
                     19703 => "00100101",
                     19704 => "00100111",
                     19705 => "00101000",
                     19706 => "00000000",
                     19707 => "00001001",
                     19708 => "00010010",
                     19709 => "00011011",
                     19710 => "00100001",
                     19711 => "00100111",
                     19712 => "00101100",
                     19713 => "00101111",
                     19714 => "00110000",
                     19715 => "00000000",
                     19716 => "00001011",
                     19717 => "00010101",
                     19718 => "00011111",
                     19719 => "00100111",
                     19720 => "00101110",
                     19721 => "00110011",
                     19722 => "00110111",
                     19723 => "00111000",
                     19724 => "00000000",
                     19725 => "00001100",
                     19726 => "00011000",
                     19727 => "00100100",
                     19728 => "00101101",
                     19729 => "00110101",
                     19730 => "00111011",
                     19731 => "00111110",
                     19732 => "01000000",
                     19733 => "00000000",
                     19734 => "00001110",
                     19735 => "00011011",
                     19736 => "00101000",
                     19737 => "00110010",
                     19738 => "00111011",
                     19739 => "01000010",
                     19740 => "01000110",
                     19741 => "01001000",
                     19742 => "00000000",
                     19743 => "00001111",
                     19744 => "00011111",
                     19745 => "00101101",
                     19746 => "00111000",
                     19747 => "01000010",
                     19748 => "01001010",
                     19749 => "01001110",
                     19750 => "01010000",
                     19751 => "00000000",
                     19752 => "00010001",
                     19753 => "00100010",
                     19754 => "00110001",
                     19755 => "00111110",
                     19756 => "01001001",
                     19757 => "01010001",
                     19758 => "01010110",
                     19759 => "01011000",
                     19760 => "00000001",
                     19761 => "00000011",
                     19762 => "00000010",
                     19763 => "00000000",
                     19764 => "00000000",
                     19765 => "00001001",
                     19766 => "00010010",
                     19767 => "00011011",
                     19768 => "00100100",
                     19769 => "00101101",
                     19770 => "00110110",
                     19771 => "00111111",
                     19772 => "01001000",
                     19773 => "01010001",
                     19774 => "01011010",
                     19775 => "01100011",
                     19776 => "00001100",
                     19777 => "00011000",
                     19778 => "00100000",
                     19779 => "10110110",
                     19780 => "11110001",
                     19781 => "10101101",
                     19782 => "11010001",
                     19783 => "00000011",
                     19784 => "00101001",
                     19785 => "00001000",
                     19786 => "11010000",
                     19787 => "01110100",
                     19788 => "10101101",
                     19789 => "01000111",
                     19790 => "00000111",
                     19791 => "11010000",
                     19792 => "00001010",
                     19793 => "10111101",
                     19794 => "10001000",
                     19795 => "00000011",
                     19796 => "00100000",
                     19797 => "11011000",
                     19798 => "11010011",
                     19799 => "00101001",
                     19800 => "00011111",
                     19801 => "10010101",
                     19802 => "10100000",
                     19803 => "10110101",
                     19804 => "10100000",
                     19805 => "10110100",
                     19806 => "00010110",
                     19807 => "11000000",
                     19808 => "00011111",
                     19809 => "10010000",
                     19810 => "00001101",
                     19811 => "11001001",
                     19812 => "00001000",
                     19813 => "11110000",
                     19814 => "00000100",
                     19815 => "11001001",
                     19816 => "00011000",
                     19817 => "11010000",
                     19818 => "00000101",
                     19819 => "00011000",
                     19820 => "01101001",
                     19821 => "00000001",
                     19822 => "10010101",
                     19823 => "10100000",
                     19824 => "10000101",
                     19825 => "11101111",
                     19826 => "00100000",
                     19827 => "01011001",
                     19828 => "11110001",
                     19829 => "00100000",
                     19830 => "10010100",
                     19831 => "11001110",
                     19832 => "10111100",
                     19833 => "11100101",
                     19834 => "00000110",
                     19835 => "10101101",
                     19836 => "10111001",
                     19837 => "00000011",
                     19838 => "10011001",
                     19839 => "00000000",
                     19840 => "00000010",
                     19841 => "10000101",
                     19842 => "00000111",
                     19843 => "10101101",
                     19844 => "10101110",
                     19845 => "00000011",
                     19846 => "10011001",
                     19847 => "00000011",
                     19848 => "00000010",
                     19849 => "10000101",
                     19850 => "00000110",
                     19851 => "10101001",
                     19852 => "00000001",
                     19853 => "10000101",
                     19854 => "00000000",
                     19855 => "00100000",
                     19856 => "00001110",
                     19857 => "11001110",
                     19858 => "10100000",
                     19859 => "00000101",
                     19860 => "10110101",
                     19861 => "00010110",
                     19862 => "11001001",
                     19863 => "00011111",
                     19864 => "10010000",
                     19865 => "00000010",
                     19866 => "10100000",
                     19867 => "00001011",
                     19868 => "10000100",
                     19869 => "11101101",
                     19870 => "10101001",
                     19871 => "00000000",
                     19872 => "10000101",
                     19873 => "00000000",
                     19874 => "10100101",
                     19875 => "11101111",
                     19876 => "00100000",
                     19877 => "10010100",
                     19878 => "11001110",
                     19879 => "00100000",
                     19880 => "11000001",
                     19881 => "11001101",
                     19882 => "10100101",
                     19883 => "00000000",
                     19884 => "11001001",
                     19885 => "00000100",
                     19886 => "11010000",
                     19887 => "00001000",
                     19888 => "10101100",
                     19889 => "11001111",
                     19890 => "00000110",
                     19891 => "10111001",
                     19892 => "11100101",
                     19893 => "00000110",
                     19894 => "10000101",
                     19895 => "00000110",
                     19896 => "11100110",
                     19897 => "00000000",
                     19898 => "10100101",
                     19899 => "00000000",
                     19900 => "11000101",
                     19901 => "11101101",
                     19902 => "10010000",
                     19903 => "11100010",
                     19904 => "01100000",
                     19905 => "10100101",
                     19906 => "00000011",
                     19907 => "10000101",
                     19908 => "00000101",
                     19909 => "10100100",
                     19910 => "00000110",
                     19911 => "10100101",
                     19912 => "00000001",
                     19913 => "01000110",
                     19914 => "00000101",
                     19915 => "10110000",
                     19916 => "00000100",
                     19917 => "01001001",
                     19918 => "11111111",
                     19919 => "01101001",
                     19920 => "00000001",
                     19921 => "00011000",
                     19922 => "01101101",
                     19923 => "10101110",
                     19924 => "00000011",
                     19925 => "10011001",
                     19926 => "00000011",
                     19927 => "00000010",
                     19928 => "10000101",
                     19929 => "00000110",
                     19930 => "11001101",
                     19931 => "10101110",
                     19932 => "00000011",
                     19933 => "10110000",
                     19934 => "00001001",
                     19935 => "10101101",
                     19936 => "10101110",
                     19937 => "00000011",
                     19938 => "00111000",
                     19939 => "11100101",
                     19940 => "00000110",
                     19941 => "01001100",
                     19942 => "11101100",
                     19943 => "11001101",
                     19944 => "00111000",
                     19945 => "11101101",
                     19946 => "10101110",
                     19947 => "00000011",
                     19948 => "11001001",
                     19949 => "01011001",
                     19950 => "10010000",
                     19951 => "00000100",
                     19952 => "10101001",
                     19953 => "11111000",
                     19954 => "11010000",
                     19955 => "00010101",
                     19956 => "10101101",
                     19957 => "10111001",
                     19958 => "00000011",
                     19959 => "11001001",
                     19960 => "11111000",
                     19961 => "11110000",
                     19962 => "00001110",
                     19963 => "10100101",
                     19964 => "00000010",
                     19965 => "01000110",
                     19966 => "00000101",
                     19967 => "10110000",
                     19968 => "00000100",
                     19969 => "01001001",
                     19970 => "11111111",
                     19971 => "01101001",
                     19972 => "00000001",
                     19973 => "00011000",
                     19974 => "01101101",
                     19975 => "10111001",
                     19976 => "00000011",
                     19977 => "10011001",
                     19978 => "00000000",
                     19979 => "00000010",
                     19980 => "10000101",
                     19981 => "00000111",
                     19982 => "00100000",
                     19983 => "11110100",
                     19984 => "11101100",
                     19985 => "10011000",
                     19986 => "01001000",
                     19987 => "10101101",
                     19988 => "10011111",
                     19989 => "00000111",
                     19990 => "00001101",
                     19991 => "01000111",
                     19992 => "00000111",
                     19993 => "11010000",
                     19994 => "01110000",
                     19995 => "10000101",
                     19996 => "00000101",
                     19997 => "10100100",
                     19998 => "10110101",
                     19999 => "10001000",
                     20000 => "11010000",
                     20001 => "01101001",
                     20002 => "10100100",
                     20003 => "11001110",
                     20004 => "10101101",
                     20005 => "01010100",
                     20006 => "00000111",
                     20007 => "11010000",
                     20008 => "00000101",
                     20009 => "10101101",
                     20010 => "00010100",
                     20011 => "00000111",
                     20012 => "11110000",
                     20013 => "00001001",
                     20014 => "11100110",
                     20015 => "00000101",
                     20016 => "11100110",
                     20017 => "00000101",
                     20018 => "10011000",
                     20019 => "00011000",
                     20020 => "01101001",
                     20021 => "00011000",
                     20022 => "10101000",
                     20023 => "10011000",
                     20024 => "00111000",
                     20025 => "11100101",
                     20026 => "00000111",
                     20027 => "00010000",
                     20028 => "00000101",
                     20029 => "01001001",
                     20030 => "11111111",
                     20031 => "00011000",
                     20032 => "01101001",
                     20033 => "00000001",
                     20034 => "11001001",
                     20035 => "00001000",
                     20036 => "10110000",
                     20037 => "00011100",
                     20038 => "10100101",
                     20039 => "00000110",
                     20040 => "11001001",
                     20041 => "11110000",
                     20042 => "10110000",
                     20043 => "00010110",
                     20044 => "10101101",
                     20045 => "00000111",
                     20046 => "00000010",
                     20047 => "00011000",
                     20048 => "01101001",
                     20049 => "00000100",
                     20050 => "10000101",
                     20051 => "00000100",
                     20052 => "00111000",
                     20053 => "11100101",
                     20054 => "00000110",
                     20055 => "00010000",
                     20056 => "00000101",
                     20057 => "01001001",
                     20058 => "11111111",
                     20059 => "00011000",
                     20060 => "01101001",
                     20061 => "00000001",
                     20062 => "11001001",
                     20063 => "00001000",
                     20064 => "10010000",
                     20065 => "00010011",
                     20066 => "10100101",
                     20067 => "00000101",
                     20068 => "11001001",
                     20069 => "00000010",
                     20070 => "11110000",
                     20071 => "00100011",
                     20072 => "10100100",
                     20073 => "00000101",
                     20074 => "10100101",
                     20075 => "11001110",
                     20076 => "00011000",
                     20077 => "01111001",
                     20078 => "01000000",
                     20079 => "11001101",
                     20080 => "11100110",
                     20081 => "00000101",
                     20082 => "01001100",
                     20083 => "00111000",
                     20084 => "11001110",
                     20085 => "10100010",
                     20086 => "00000001",
                     20087 => "10100101",
                     20088 => "00000100",
                     20089 => "11000101",
                     20090 => "00000110",
                     20091 => "10110000",
                     20092 => "00000001",
                     20093 => "11101000",
                     20094 => "10000110",
                     20095 => "01000110",
                     20096 => "10100010",
                     20097 => "00000000",
                     20098 => "10100101",
                     20099 => "00000000",
                     20100 => "01001000",
                     20101 => "00100000",
                     20102 => "00101101",
                     20103 => "11011001",
                     20104 => "01101000",
                     20105 => "10000101",
                     20106 => "00000000",
                     20107 => "01101000",
                     20108 => "00011000",
                     20109 => "01101001",
                     20110 => "00000100",
                     20111 => "10000101",
                     20112 => "00000110",
                     20113 => "10100110",
                     20114 => "00001000",
                     20115 => "01100000",
                     20116 => "01001000",
                     20117 => "00101001",
                     20118 => "00001111",
                     20119 => "11001001",
                     20120 => "00001001",
                     20121 => "10010000",
                     20122 => "00000101",
                     20123 => "01001001",
                     20124 => "00001111",
                     20125 => "00011000",
                     20126 => "01101001",
                     20127 => "00000001",
                     20128 => "10000101",
                     20129 => "00000001",
                     20130 => "10100100",
                     20131 => "00000000",
                     20132 => "10111001",
                     20133 => "00110100",
                     20134 => "11001101",
                     20135 => "00011000",
                     20136 => "01100101",
                     20137 => "00000001",
                     20138 => "10101000",
                     20139 => "10111001",
                     20140 => "11001101",
                     20141 => "11001100",
                     20142 => "10000101",
                     20143 => "00000001",
                     20144 => "01101000",
                     20145 => "01001000",
                     20146 => "00011000",
                     20147 => "01101001",
                     20148 => "00001000",
                     20149 => "00101001",
                     20150 => "00001111",
                     20151 => "11001001",
                     20152 => "00001001",
                     20153 => "10010000",
                     20154 => "00000101",
                     20155 => "01001001",
                     20156 => "00001111",
                     20157 => "00011000",
                     20158 => "01101001",
                     20159 => "00000001",
                     20160 => "10000101",
                     20161 => "00000010",
                     20162 => "10100100",
                     20163 => "00000000",
                     20164 => "10111001",
                     20165 => "00110100",
                     20166 => "11001101",
                     20167 => "00011000",
                     20168 => "01100101",
                     20169 => "00000010",
                     20170 => "10101000",
                     20171 => "10111001",
                     20172 => "11001101",
                     20173 => "11001100",
                     20174 => "10000101",
                     20175 => "00000010",
                     20176 => "01101000",
                     20177 => "01001010",
                     20178 => "01001010",
                     20179 => "01001010",
                     20180 => "10101000",
                     20181 => "10111001",
                     20182 => "00110000",
                     20183 => "11001101",
                     20184 => "10000101",
                     20185 => "00000011",
                     20186 => "01100000",
                     20187 => "10100000",
                     20188 => "00100000",
                     20189 => "10110101",
                     20190 => "00011110",
                     20191 => "00101001",
                     20192 => "00100000",
                     20193 => "11010000",
                     20194 => "00000101",
                     20195 => "00100000",
                     20196 => "00000111",
                     20197 => "10111111",
                     20198 => "10100000",
                     20199 => "00010111",
                     20200 => "10101001",
                     20201 => "00000101",
                     20202 => "01001100",
                     20203 => "10011011",
                     20204 => "10111111",
                     20205 => "00010101",
                     20206 => "00110000",
                     20207 => "01000000",
                     20208 => "10110101",
                     20209 => "00011110",
                     20210 => "00101001",
                     20211 => "00100000",
                     20212 => "11110000",
                     20213 => "00000011",
                     20214 => "01001100",
                     20215 => "01101000",
                     20216 => "10111111",
                     20217 => "10110101",
                     20218 => "00011110",
                     20219 => "11110000",
                     20220 => "00001011",
                     20221 => "10101001",
                     20222 => "00000000",
                     20223 => "10010101",
                     20224 => "10100000",
                     20225 => "10001101",
                     20226 => "11001011",
                     20227 => "00000110",
                     20228 => "10101001",
                     20229 => "00010000",
                     20230 => "11010000",
                     20231 => "00010011",
                     20232 => "10101001",
                     20233 => "00010010",
                     20234 => "10001101",
                     20235 => "11001011",
                     20236 => "00000110",
                     20237 => "10100000",
                     20238 => "00000010",
                     20239 => "10111001",
                     20240 => "11101101",
                     20241 => "11001110",
                     20242 => "10011001",
                     20243 => "00000001",
                     20244 => "00000000",
                     20245 => "10001000",
                     20246 => "00010000",
                     20247 => "11110111",
                     20248 => "00100000",
                     20249 => "00110100",
                     20250 => "11001111",
                     20251 => "10010101",
                     20252 => "01011000",
                     20253 => "10100000",
                     20254 => "00000001",
                     20255 => "10110101",
                     20256 => "10100000",
                     20257 => "00101001",
                     20258 => "00000001",
                     20259 => "11010000",
                     20260 => "00001010",
                     20261 => "10110101",
                     20262 => "01011000",
                     20263 => "01001001",
                     20264 => "11111111",
                     20265 => "00011000",
                     20266 => "01101001",
                     20267 => "00000001",
                     20268 => "10010101",
                     20269 => "01011000",
                     20270 => "11001000",
                     20271 => "10010100",
                     20272 => "01000110",
                     20273 => "01001100",
                     20274 => "00000111",
                     20275 => "10111111",
                     20276 => "10100000",
                     20277 => "00000000",
                     20278 => "00100000",
                     20279 => "01001011",
                     20280 => "11100001",
                     20281 => "00010000",
                     20282 => "00001010",
                     20283 => "11001000",
                     20284 => "10100101",
                     20285 => "00000000",
                     20286 => "01001001",
                     20287 => "11111111",
                     20288 => "00011000",
                     20289 => "01101001",
                     20290 => "00000001",
                     20291 => "10000101",
                     20292 => "00000000",
                     20293 => "10100101",
                     20294 => "00000000",
                     20295 => "11001001",
                     20296 => "00111100",
                     20297 => "10010000",
                     20298 => "00011100",
                     20299 => "10101001",
                     20300 => "00111100",
                     20301 => "10000101",
                     20302 => "00000000",
                     20303 => "10110101",
                     20304 => "00010110",
                     20305 => "11001001",
                     20306 => "00010001",
                     20307 => "11010000",
                     20308 => "00010010",
                     20309 => "10011000",
                     20310 => "11010101",
                     20311 => "10100000",
                     20312 => "11110000",
                     20313 => "00001101",
                     20314 => "10110101",
                     20315 => "10100000",
                     20316 => "11110000",
                     20317 => "00000110",
                     20318 => "11010110",
                     20319 => "01011000",
                     20320 => "10110101",
                     20321 => "01011000",
                     20322 => "11010000",
                     20323 => "01000000",
                     20324 => "10011000",
                     20325 => "10010101",
                     20326 => "10100000",
                     20327 => "10100101",
                     20328 => "00000000",
                     20329 => "00101001",
                     20330 => "00111100",
                     20331 => "01001010",
                     20332 => "01001010",
                     20333 => "10000101",
                     20334 => "00000000",
                     20335 => "10100000",
                     20336 => "00000000",
                     20337 => "10100101",
                     20338 => "01010111",
                     20339 => "11110000",
                     20340 => "00100100",
                     20341 => "10101101",
                     20342 => "01110101",
                     20343 => "00000111",
                     20344 => "11110000",
                     20345 => "00011111",
                     20346 => "11001000",
                     20347 => "10100101",
                     20348 => "01010111",
                     20349 => "11001001",
                     20350 => "00011101",
                     20351 => "10010000",
                     20352 => "00001000",
                     20353 => "10101101",
                     20354 => "01110101",
                     20355 => "00000111",
                     20356 => "11001001",
                     20357 => "00000010",
                     20358 => "10010000",
                     20359 => "00000001",
                     20360 => "11001000",
                     20361 => "10110101",
                     20362 => "00010110",
                     20363 => "11001001",
                     20364 => "00010010",
                     20365 => "11010000",
                     20366 => "00000100",
                     20367 => "10100101",
                     20368 => "01010111",
                     20369 => "11010000",
                     20370 => "00000110",
                     20371 => "10110101",
                     20372 => "10100000",
                     20373 => "11010000",
                     20374 => "00000010",
                     20375 => "10100000",
                     20376 => "00000000",
                     20377 => "10111001",
                     20378 => "00000001",
                     20379 => "00000000",
                     20380 => "10100100",
                     20381 => "00000000",
                     20382 => "00111000",
                     20383 => "11101001",
                     20384 => "00000001",
                     20385 => "10001000",
                     20386 => "00010000",
                     20387 => "11111010",
                     20388 => "01100000",
                     20389 => "00011010",
                     20390 => "01011000",
                     20391 => "10011000",
                     20392 => "10010110",
                     20393 => "10010100",
                     20394 => "10010010",
                     20395 => "10010000",
                     20396 => "10001110",
                     20397 => "10001100",
                     20398 => "10001010",
                     20399 => "10001000",
                     20400 => "10000110",
                     20401 => "10000100",
                     20402 => "10000010",
                     20403 => "10000000",
                     20404 => "10101110",
                     20405 => "01101000",
                     20406 => "00000011",
                     20407 => "10110101",
                     20408 => "00010110",
                     20409 => "11001001",
                     20410 => "00101101",
                     20411 => "11010000",
                     20412 => "00010000",
                     20413 => "10000110",
                     20414 => "00001000",
                     20415 => "10110101",
                     20416 => "00011110",
                     20417 => "11110000",
                     20418 => "00011010",
                     20419 => "00101001",
                     20420 => "01000000",
                     20421 => "11110000",
                     20422 => "00000110",
                     20423 => "10110101",
                     20424 => "11001111",
                     20425 => "11001001",
                     20426 => "11100000",
                     20427 => "10010000",
                     20428 => "00001010",
                     20429 => "10101001",
                     20430 => "10000000",
                     20431 => "10000101",
                     20432 => "11111100",
                     20433 => "11101110",
                     20434 => "01110010",
                     20435 => "00000111",
                     20436 => "01001100",
                     20437 => "00111001",
                     20438 => "11010000",
                     20439 => "00100000",
                     20440 => "10010001",
                     20441 => "10111111",
                     20442 => "01001100",
                     20443 => "01000011",
                     20444 => "11010001",
                     20445 => "11001110",
                     20446 => "01100100",
                     20447 => "00000011",
                     20448 => "11010000",
                     20449 => "01000100",
                     20450 => "10101001",
                     20451 => "00000100",
                     20452 => "10001101",
                     20453 => "01100100",
                     20454 => "00000011",
                     20455 => "10101101",
                     20456 => "01100011",
                     20457 => "00000011",
                     20458 => "01001001",
                     20459 => "00000001",
                     20460 => "10001101",
                     20461 => "01100011",
                     20462 => "00000011",
                     20463 => "10101001",
                     20464 => "00100010",
                     20465 => "10000101",
                     20466 => "00000101",
                     20467 => "10101100",
                     20468 => "01101001",
                     20469 => "00000011",
                     20470 => "10111001",
                     20471 => "10100101",
                     20472 => "11001111",
                     20473 => "10000101",
                     20474 => "00000100",
                     20475 => "10101100",
                     20476 => "00000000",
                     20477 => "00000011",
                     20478 => "11001000",
                     20479 => "10100010",
                     20480 => "00001100",
                     20481 => "00100000",
                     20482 => "11001101",
                     20483 => "10001010",
                     20484 => "10100110",
                     20485 => "00001000",
                     20486 => "00100000",
                     20487 => "10001111",
                     20488 => "10001010",
                     20489 => "10101001",
                     20490 => "00001000",
                     20491 => "10000101",
                     20492 => "11111110",
                     20493 => "10101001",
                     20494 => "00000001",
                     20495 => "10000101",
                     20496 => "11111101",
                     20497 => "11101110",
                     20498 => "01101001",
                     20499 => "00000011",
                     20500 => "10101101",
                     20501 => "01101001",
                     20502 => "00000011",
                     20503 => "11001001",
                     20504 => "00001111",
                     20505 => "11010000",
                     20506 => "00001011",
                     20507 => "00100000",
                     20508 => "01101001",
                     20509 => "11000011",
                     20510 => "10101001",
                     20511 => "01000000",
                     20512 => "10010101",
                     20513 => "00011110",
                     20514 => "10101001",
                     20515 => "10000000",
                     20516 => "10000101",
                     20517 => "11111110",
                     20518 => "01001100",
                     20519 => "01000011",
                     20520 => "11010001",
                     20521 => "00100001",
                     20522 => "01000001",
                     20523 => "00010001",
                     20524 => "00110001",
                     20525 => "10110101",
                     20526 => "00011110",
                     20527 => "00101001",
                     20528 => "00100000",
                     20529 => "11110000",
                     20530 => "00010100",
                     20531 => "10110101",
                     20532 => "11001111",
                     20533 => "11001001",
                     20534 => "11100000",
                     20535 => "10010000",
                     20536 => "10011110",
                     20537 => "10100010",
                     20538 => "00000100",
                     20539 => "00100000",
                     20540 => "10011110",
                     20541 => "11001001",
                     20542 => "11001010",
                     20543 => "00010000",
                     20544 => "11111010",
                     20545 => "10001101",
                     20546 => "11001011",
                     20547 => "00000110",
                     20548 => "10100110",
                     20549 => "00001000",
                     20550 => "01100000",
                     20551 => "10101001",
                     20552 => "00000000",
                     20553 => "10001101",
                     20554 => "11001011",
                     20555 => "00000110",
                     20556 => "10101101",
                     20557 => "01000111",
                     20558 => "00000111",
                     20559 => "11110000",
                     20560 => "00000011",
                     20561 => "01001100",
                     20562 => "00000001",
                     20563 => "11010001",
                     20564 => "10101101",
                     20565 => "01100011",
                     20566 => "00000011",
                     20567 => "00010000",
                     20568 => "00000011",
                     20569 => "01001100",
                     20570 => "11010111",
                     20571 => "11010000",
                     20572 => "11001110",
                     20573 => "01100100",
                     20574 => "00000011",
                     20575 => "11010000",
                     20576 => "00001101",
                     20577 => "10101001",
                     20578 => "00100000",
                     20579 => "10001101",
                     20580 => "01100100",
                     20581 => "00000011",
                     20582 => "10101101",
                     20583 => "01100011",
                     20584 => "00000011",
                     20585 => "01001001",
                     20586 => "00000001",
                     20587 => "10001101",
                     20588 => "01100011",
                     20589 => "00000011",
                     20590 => "10100101",
                     20591 => "00001001",
                     20592 => "00101001",
                     20593 => "00001111",
                     20594 => "11010000",
                     20595 => "00000100",
                     20596 => "10101001",
                     20597 => "00000010",
                     20598 => "10010101",
                     20599 => "01000110",
                     20600 => "10111101",
                     20601 => "10001010",
                     20602 => "00000111",
                     20603 => "11110000",
                     20604 => "00011100",
                     20605 => "00100000",
                     20606 => "01001011",
                     20607 => "11100001",
                     20608 => "00010000",
                     20609 => "00010111",
                     20610 => "10101001",
                     20611 => "00000001",
                     20612 => "10010101",
                     20613 => "01000110",
                     20614 => "10101001",
                     20615 => "00000010",
                     20616 => "10001101",
                     20617 => "01100101",
                     20618 => "00000011",
                     20619 => "10101001",
                     20620 => "00100000",
                     20621 => "10011101",
                     20622 => "10001010",
                     20623 => "00000111",
                     20624 => "10001101",
                     20625 => "10010000",
                     20626 => "00000111",
                     20627 => "10110101",
                     20628 => "10000111",
                     20629 => "11001001",
                     20630 => "11001000",
                     20631 => "10110000",
                     20632 => "00111110",
                     20633 => "10100101",
                     20634 => "00001001",
                     20635 => "00101001",
                     20636 => "00000011",
                     20637 => "11010000",
                     20638 => "00111000",
                     20639 => "10110101",
                     20640 => "10000111",
                     20641 => "11001101",
                     20642 => "01100110",
                     20643 => "00000011",
                     20644 => "11010000",
                     20645 => "00001100",
                     20646 => "10111101",
                     20647 => "10100111",
                     20648 => "00000111",
                     20649 => "00101001",
                     20650 => "00000011",
                     20651 => "10101000",
                     20652 => "10111001",
                     20653 => "00101001",
                     20654 => "11010000",
                     20655 => "10001101",
                     20656 => "11011100",
                     20657 => "00000110",
                     20658 => "10110101",
                     20659 => "10000111",
                     20660 => "00011000",
                     20661 => "01101101",
                     20662 => "01100101",
                     20663 => "00000011",
                     20664 => "10010101",
                     20665 => "10000111",
                     20666 => "10110100",
                     20667 => "01000110",
                     20668 => "11000000",
                     20669 => "00000001",
                     20670 => "11110000",
                     20671 => "00010111",
                     20672 => "10100000",
                     20673 => "11111111",
                     20674 => "00111000",
                     20675 => "11101101",
                     20676 => "01100110",
                     20677 => "00000011",
                     20678 => "00010000",
                     20679 => "00000111",
                     20680 => "01001001",
                     20681 => "11111111",
                     20682 => "00011000",
                     20683 => "01101001",
                     20684 => "00000001",
                     20685 => "10100000",
                     20686 => "00000001",
                     20687 => "11001101",
                     20688 => "11011100",
                     20689 => "00000110",
                     20690 => "10010000",
                     20691 => "00000011",
                     20692 => "10001100",
                     20693 => "01100101",
                     20694 => "00000011",
                     20695 => "10111101",
                     20696 => "10001010",
                     20697 => "00000111",
                     20698 => "11010000",
                     20699 => "00101000",
                     20700 => "00100000",
                     20701 => "10010001",
                     20702 => "10111111",
                     20703 => "10101101",
                     20704 => "01011111",
                     20705 => "00000111",
                     20706 => "11001001",
                     20707 => "00000101",
                     20708 => "10010000",
                     20709 => "00001001",
                     20710 => "10100101",
                     20711 => "00001001",
                     20712 => "00101001",
                     20713 => "00000011",
                     20714 => "11010000",
                     20715 => "00000011",
                     20716 => "00100000",
                     20717 => "10011001",
                     20718 => "10111010",
                     20719 => "10110101",
                     20720 => "11001111",
                     20721 => "11001001",
                     20722 => "10000000",
                     20723 => "10010000",
                     20724 => "00011100",
                     20725 => "10111101",
                     20726 => "10100111",
                     20727 => "00000111",
                     20728 => "00101001",
                     20729 => "00000011",
                     20730 => "10101000",
                     20731 => "10111001",
                     20732 => "00101001",
                     20733 => "11010000",
                     20734 => "10011101",
                     20735 => "10001010",
                     20736 => "00000111",
                     20737 => "01001100",
                     20738 => "00010001",
                     20739 => "11010001",
                     20740 => "11001001",
                     20741 => "00000001",
                     20742 => "11010000",
                     20743 => "00001001",
                     20744 => "11010110",
                     20745 => "11001111",
                     20746 => "00100000",
                     20747 => "01101001",
                     20748 => "11000011",
                     20749 => "10101001",
                     20750 => "11111110",
                     20751 => "10010101",
                     20752 => "10100000",
                     20753 => "10101101",
                     20754 => "01011111",
                     20755 => "00000111",
                     20756 => "11001001",
                     20757 => "00000111",
                     20758 => "11110000",
                     20759 => "00000100",
                     20760 => "11001001",
                     20761 => "00000101",
                     20762 => "10110000",
                     20763 => "00100111",
                     20764 => "10101101",
                     20765 => "10010000",
                     20766 => "00000111",
                     20767 => "11010000",
                     20768 => "00100010",
                     20769 => "10101001",
                     20770 => "00100000",
                     20771 => "10001101",
                     20772 => "10010000",
                     20773 => "00000111",
                     20774 => "10101101",
                     20775 => "01100011",
                     20776 => "00000011",
                     20777 => "01001001",
                     20778 => "10000000",
                     20779 => "10001101",
                     20780 => "01100011",
                     20781 => "00000011",
                     20782 => "00110000",
                     20783 => "11100001",
                     20784 => "00100000",
                     20785 => "10100001",
                     20786 => "11010001",
                     20787 => "10101100",
                     20788 => "11001100",
                     20789 => "00000110",
                     20790 => "11110000",
                     20791 => "00000011",
                     20792 => "00111000",
                     20793 => "11101001",
                     20794 => "00010000",
                     20795 => "10001101",
                     20796 => "10010000",
                     20797 => "00000111",
                     20798 => "10101001",
                     20799 => "00010101",
                     20800 => "10001101",
                     20801 => "11001011",
                     20802 => "00000110",
                     20803 => "00100000",
                     20804 => "10000100",
                     20805 => "11010001",
                     20806 => "10100000",
                     20807 => "00010000",
                     20808 => "10110101",
                     20809 => "01000110",
                     20810 => "01001010",
                     20811 => "10010000",
                     20812 => "00000010",
                     20813 => "10100000",
                     20814 => "11110000",
                     20815 => "10011000",
                     20816 => "00011000",
                     20817 => "01110101",
                     20818 => "10000111",
                     20819 => "10101100",
                     20820 => "11001111",
                     20821 => "00000110",
                     20822 => "10011001",
                     20823 => "10000111",
                     20824 => "00000000",
                     20825 => "10110101",
                     20826 => "11001111",
                     20827 => "00011000",
                     20828 => "01101001",
                     20829 => "00001000",
                     20830 => "10011001",
                     20831 => "11001111",
                     20832 => "00000000",
                     20833 => "10110101",
                     20834 => "00011110",
                     20835 => "10011001",
                     20836 => "00011110",
                     20837 => "00000000",
                     20838 => "10110101",
                     20839 => "01000110",
                     20840 => "10011001",
                     20841 => "01000110",
                     20842 => "00000000",
                     20843 => "10100101",
                     20844 => "00001000",
                     20845 => "01001000",
                     20846 => "10101110",
                     20847 => "11001111",
                     20848 => "00000110",
                     20849 => "10000110",
                     20850 => "00001000",
                     20851 => "10101001",
                     20852 => "00101101",
                     20853 => "10010101",
                     20854 => "00010110",
                     20855 => "00100000",
                     20856 => "10000100",
                     20857 => "11010001",
                     20858 => "01101000",
                     20859 => "10000101",
                     20860 => "00001000",
                     20861 => "10101010",
                     20862 => "10101001",
                     20863 => "00000000",
                     20864 => "10001101",
                     20865 => "01101010",
                     20866 => "00000011",
                     20867 => "01100000",
                     20868 => "11101110",
                     20869 => "01101010",
                     20870 => "00000011",
                     20871 => "00100000",
                     20872 => "11011101",
                     20873 => "11001000",
                     20874 => "10110101",
                     20875 => "00011110",
                     20876 => "11010000",
                     20877 => "11110101",
                     20878 => "10101001",
                     20879 => "00001010",
                     20880 => "10011101",
                     20881 => "10011010",
                     20882 => "00000100",
                     20883 => "00100000",
                     20884 => "01001011",
                     20885 => "11100010",
                     20886 => "01001100",
                     20887 => "01010011",
                     20888 => "11011000",
                     20889 => "10000000",
                     20890 => "00110000",
                     20891 => "00110000",
                     20892 => "10000000",
                     20893 => "10000000",
                     20894 => "10000000",
                     20895 => "00110000",
                     20896 => "01010000",
                     20897 => "10101100",
                     20898 => "01100111",
                     20899 => "00000011",
                     20900 => "11101110",
                     20901 => "01100111",
                     20902 => "00000011",
                     20903 => "10101101",
                     20904 => "01100111",
                     20905 => "00000011",
                     20906 => "00101001",
                     20907 => "00000111",
                     20908 => "10001101",
                     20909 => "01100111",
                     20910 => "00000011",
                     20911 => "10111001",
                     20912 => "10011001",
                     20913 => "11010001",
                     20914 => "01100000",
                     20915 => "10101101",
                     20916 => "01000111",
                     20917 => "00000111",
                     20918 => "11010000",
                     20919 => "00110000",
                     20920 => "10101001",
                     20921 => "01110000",
                     20922 => "10101100",
                     20923 => "11001100",
                     20924 => "00000110",
                     20925 => "11110000",
                     20926 => "00000010",
                     20927 => "10101001",
                     20928 => "10010000",
                     20929 => "10000101",
                     20930 => "00000000",
                     20931 => "10111101",
                     20932 => "00000001",
                     20933 => "00000100",
                     20934 => "00111000",
                     20935 => "11100101",
                     20936 => "00000000",
                     20937 => "10011101",
                     20938 => "00000001",
                     20939 => "00000100",
                     20940 => "10110101",
                     20941 => "10000111",
                     20942 => "11101001",
                     20943 => "00000001",
                     20944 => "10010101",
                     20945 => "10000111",
                     20946 => "10110101",
                     20947 => "01101110",
                     20948 => "11101001",
                     20949 => "00000000",
                     20950 => "10010101",
                     20951 => "01101110",
                     20952 => "10111100",
                     20953 => "00010111",
                     20954 => "00000100",
                     20955 => "10110101",
                     20956 => "11001111",
                     20957 => "11011001",
                     20958 => "10100011",
                     20959 => "11000101",
                     20960 => "11110000",
                     20961 => "00000110",
                     20962 => "00011000",
                     20963 => "01111101",
                     20964 => "00110100",
                     20965 => "00000100",
                     20966 => "10010101",
                     20967 => "11001111",
                     20968 => "00100000",
                     20969 => "01011001",
                     20970 => "11110001",
                     20971 => "10110101",
                     20972 => "00011110",
                     20973 => "11010000",
                     20974 => "11000011",
                     20975 => "10101001",
                     20976 => "01010001",
                     20977 => "10000101",
                     20978 => "00000000",
                     20979 => "10100000",
                     20980 => "00000010",
                     20981 => "10100101",
                     20982 => "00001001",
                     20983 => "00101001",
                     20984 => "00000010",
                     20985 => "11110000",
                     20986 => "00000010",
                     20987 => "10100000",
                     20988 => "10000010",
                     20989 => "10000100",
                     20990 => "00000001",
                     20991 => "10111100",
                     20992 => "11100101",
                     20993 => "00000110",
                     20994 => "10100010",
                     20995 => "00000000",
                     20996 => "10101101",
                     20997 => "10111001",
                     20998 => "00000011",
                     20999 => "10011001",
                     21000 => "00000000",
                     21001 => "00000010",
                     21002 => "10100101",
                     21003 => "00000000",
                     21004 => "10011001",
                     21005 => "00000001",
                     21006 => "00000010",
                     21007 => "11100110",
                     21008 => "00000000",
                     21009 => "10100101",
                     21010 => "00000001",
                     21011 => "10011001",
                     21012 => "00000010",
                     21013 => "00000010",
                     21014 => "10101101",
                     21015 => "10101110",
                     21016 => "00000011",
                     21017 => "10011001",
                     21018 => "00000011",
                     21019 => "00000010",
                     21020 => "00011000",
                     21021 => "01101001",
                     21022 => "00001000",
                     21023 => "10001101",
                     21024 => "10101110",
                     21025 => "00000011",
                     21026 => "11001000",
                     21027 => "11001000",
                     21028 => "11001000",
                     21029 => "11001000",
                     21030 => "11101000",
                     21031 => "11100000",
                     21032 => "00000011",
                     21033 => "10010000",
                     21034 => "11011001",
                     21035 => "10100110",
                     21036 => "00001000",
                     21037 => "00100000",
                     21038 => "10110110",
                     21039 => "11110001",
                     21040 => "10111100",
                     21041 => "11100101",
                     21042 => "00000110",
                     21043 => "10101101",
                     21044 => "11010001",
                     21045 => "00000011",
                     21046 => "01001010",
                     21047 => "01001000",
                     21048 => "10010000",
                     21049 => "00000101",
                     21050 => "10101001",
                     21051 => "11111000",
                     21052 => "10011001",
                     21053 => "00001100",
                     21054 => "00000010",
                     21055 => "01101000",
                     21056 => "01001010",
                     21057 => "01001000",
                     21058 => "10010000",
                     21059 => "00000101",
                     21060 => "10101001",
                     21061 => "11111000",
                     21062 => "10011001",
                     21063 => "00001000",
                     21064 => "00000010",
                     21065 => "01101000",
                     21066 => "01001010",
                     21067 => "01001000",
                     21068 => "10010000",
                     21069 => "00000101",
                     21070 => "10101001",
                     21071 => "11111000",
                     21072 => "10011001",
                     21073 => "00000100",
                     21074 => "00000010",
                     21075 => "01101000",
                     21076 => "01001010",
                     21077 => "10010000",
                     21078 => "00000101",
                     21079 => "10101001",
                     21080 => "11111000",
                     21081 => "10011001",
                     21082 => "00000000",
                     21083 => "00000010",
                     21084 => "01100000",
                     21085 => "11010110",
                     21086 => "10100000",
                     21087 => "11010000",
                     21088 => "00001100",
                     21089 => "10101001",
                     21090 => "00001000",
                     21091 => "10010101",
                     21092 => "10100000",
                     21093 => "11110110",
                     21094 => "01011000",
                     21095 => "10110101",
                     21096 => "01011000",
                     21097 => "11001001",
                     21098 => "00000011",
                     21099 => "10110000",
                     21100 => "00011000",
                     21101 => "00100000",
                     21102 => "01011001",
                     21103 => "11110001",
                     21104 => "10101101",
                     21105 => "10111001",
                     21106 => "00000011",
                     21107 => "10001101",
                     21108 => "10111010",
                     21109 => "00000011",
                     21110 => "10101101",
                     21111 => "10101110",
                     21112 => "00000011",
                     21113 => "10001101",
                     21114 => "10101111",
                     21115 => "00000011",
                     21116 => "10111100",
                     21117 => "11100101",
                     21118 => "00000110",
                     21119 => "10110101",
                     21120 => "01011000",
                     21121 => "00100000",
                     21122 => "00011110",
                     21123 => "11101101",
                     21124 => "01100000",
                     21125 => "10101001",
                     21126 => "00000000",
                     21127 => "10010101",
                     21128 => "00001111",
                     21129 => "10101001",
                     21130 => "00001000",
                     21131 => "10000101",
                     21132 => "11111110",
                     21133 => "10101001",
                     21134 => "00000101",
                     21135 => "10001101",
                     21136 => "00111000",
                     21137 => "00000001",
                     21138 => "01001100",
                     21139 => "11111110",
                     21140 => "11010010",
                     21141 => "00000000",
                     21142 => "00000000",
                     21143 => "00001000",
                     21144 => "00001000",
                     21145 => "00000000",
                     21146 => "00001000",
                     21147 => "00000000",
                     21148 => "00001000",
                     21149 => "01010100",
                     21150 => "01010101",
                     21151 => "01010110",
                     21152 => "01010111",
                     21153 => "10101001",
                     21154 => "00000000",
                     21155 => "10001101",
                     21156 => "11001011",
                     21157 => "00000110",
                     21158 => "10101101",
                     21159 => "01000110",
                     21160 => "00000111",
                     21161 => "11001001",
                     21162 => "00000101",
                     21163 => "10110000",
                     21164 => "00101100",
                     21165 => "00100000",
                     21166 => "00000100",
                     21167 => "10001110",
                     21168 => "11011001",
                     21169 => "11010010",
                     21170 => "10111010",
                     21171 => "11010010",
                     21172 => "11011010",
                     21173 => "11010010",
                     21174 => "00010110",
                     21175 => "11010011",
                     21176 => "01101010",
                     21177 => "11010011",
                     21178 => "10100000",
                     21179 => "00000101",
                     21180 => "10101101",
                     21181 => "11111010",
                     21182 => "00000111",
                     21183 => "11001001",
                     21184 => "00000001",
                     21185 => "11110000",
                     21186 => "00001110",
                     21187 => "10100000",
                     21188 => "00000011",
                     21189 => "11001001",
                     21190 => "00000011",
                     21191 => "11110000",
                     21192 => "00001000",
                     21193 => "10100000",
                     21194 => "00000000",
                     21195 => "11001001",
                     21196 => "00000110",
                     21197 => "11110000",
                     21198 => "00000010",
                     21199 => "10101001",
                     21200 => "11111111",
                     21201 => "10001101",
                     21202 => "11010111",
                     21203 => "00000110",
                     21204 => "10010100",
                     21205 => "00011110",
                     21206 => "11101110",
                     21207 => "01000110",
                     21208 => "00000111",
                     21209 => "01100000",
                     21210 => "10101101",
                     21211 => "11111000",
                     21212 => "00000111",
                     21213 => "00001101",
                     21214 => "11111001",
                     21215 => "00000111",
                     21216 => "00001101",
                     21217 => "11111010",
                     21218 => "00000111",
                     21219 => "11110000",
                     21220 => "11110001",
                     21221 => "10100101",
                     21222 => "00001001",
                     21223 => "00101001",
                     21224 => "00000100",
                     21225 => "11110000",
                     21226 => "00000100",
                     21227 => "10101001",
                     21228 => "00010000",
                     21229 => "10000101",
                     21230 => "11111110",
                     21231 => "10100000",
                     21232 => "00100011",
                     21233 => "10101001",
                     21234 => "11111111",
                     21235 => "10001101",
                     21236 => "00111001",
                     21237 => "00000001",
                     21238 => "00100000",
                     21239 => "01011111",
                     21240 => "10001111",
                     21241 => "10101001",
                     21242 => "00000101",
                     21243 => "10001101",
                     21244 => "00111001",
                     21245 => "00000001",
                     21246 => "10100000",
                     21247 => "00001011",
                     21248 => "10101101",
                     21249 => "01010011",
                     21250 => "00000111",
                     21251 => "11110000",
                     21252 => "00000010",
                     21253 => "10100000",
                     21254 => "00010001",
                     21255 => "00100000",
                     21256 => "01011111",
                     21257 => "10001111",
                     21258 => "10101101",
                     21259 => "01010011",
                     21260 => "00000111",
                     21261 => "00001010",
                     21262 => "00001010",
                     21263 => "00001010",
                     21264 => "00001010",
                     21265 => "00001001",
                     21266 => "00000100",
                     21267 => "01001100",
                     21268 => "00111011",
                     21269 => "10111100",
                     21270 => "10110101",
                     21271 => "11001111",
                     21272 => "11001001",
                     21273 => "01110010",
                     21274 => "10010000",
                     21275 => "00000101",
                     21276 => "11010110",
                     21277 => "11001111",
                     21278 => "01001100",
                     21279 => "00101101",
                     21280 => "11010011",
                     21281 => "10101101",
                     21282 => "11010111",
                     21283 => "00000110",
                     21284 => "11110000",
                     21285 => "00111000",
                     21286 => "00110000",
                     21287 => "00110110",
                     21288 => "10101001",
                     21289 => "00010110",
                     21290 => "10001101",
                     21291 => "11001011",
                     21292 => "00000110",
                     21293 => "00100000",
                     21294 => "01011001",
                     21295 => "11110001",
                     21296 => "10111100",
                     21297 => "11100101",
                     21298 => "00000110",
                     21299 => "10100010",
                     21300 => "00000011",
                     21301 => "10101101",
                     21302 => "10111001",
                     21303 => "00000011",
                     21304 => "00011000",
                     21305 => "01111101",
                     21306 => "10010101",
                     21307 => "11010010",
                     21308 => "10011001",
                     21309 => "00000000",
                     21310 => "00000010",
                     21311 => "10111101",
                     21312 => "10011101",
                     21313 => "11010010",
                     21314 => "10011001",
                     21315 => "00000001",
                     21316 => "00000010",
                     21317 => "10101001",
                     21318 => "00100010",
                     21319 => "10011001",
                     21320 => "00000010",
                     21321 => "00000010",
                     21322 => "10101101",
                     21323 => "10101110",
                     21324 => "00000011",
                     21325 => "00011000",
                     21326 => "01111101",
                     21327 => "10011001",
                     21328 => "11010010",
                     21329 => "10011001",
                     21330 => "00000011",
                     21331 => "00000010",
                     21332 => "11001000",
                     21333 => "11001000",
                     21334 => "11001000",
                     21335 => "11001000",
                     21336 => "11001010",
                     21337 => "00010000",
                     21338 => "11011010",
                     21339 => "10100110",
                     21340 => "00001000",
                     21341 => "01100000",
                     21342 => "00100000",
                     21343 => "00101101",
                     21344 => "11010011",
                     21345 => "10101001",
                     21346 => "00000110",
                     21347 => "10011101",
                     21348 => "10010110",
                     21349 => "00000111",
                     21350 => "11101110",
                     21351 => "01000110",
                     21352 => "00000111",
                     21353 => "01100000",
                     21354 => "00100000",
                     21355 => "00101101",
                     21356 => "11010011",
                     21357 => "10111101",
                     21358 => "10010110",
                     21359 => "00000111",
                     21360 => "11010000",
                     21361 => "00000101",
                     21362 => "10101101",
                     21363 => "10110001",
                     21364 => "00000111",
                     21365 => "11110000",
                     21366 => "11101111",
                     21367 => "01100000",
                     21368 => "10110101",
                     21369 => "00011110",
                     21370 => "11010000",
                     21371 => "01010110",
                     21372 => "10111101",
                     21373 => "10001010",
                     21374 => "00000111",
                     21375 => "11010000",
                     21376 => "01010001",
                     21377 => "10110101",
                     21378 => "10100000",
                     21379 => "11010000",
                     21380 => "00100011",
                     21381 => "10110101",
                     21382 => "01011000",
                     21383 => "00110000",
                     21384 => "00010100",
                     21385 => "00100000",
                     21386 => "01001011",
                     21387 => "11100001",
                     21388 => "00010000",
                     21389 => "00001001",
                     21390 => "10100101",
                     21391 => "00000000",
                     21392 => "01001001",
                     21393 => "11111111",
                     21394 => "00011000",
                     21395 => "01101001",
                     21396 => "00000001",
                     21397 => "10000101",
                     21398 => "00000000",
                     21399 => "10100101",
                     21400 => "00000000",
                     21401 => "11001001",
                     21402 => "00100001",
                     21403 => "10010000",
                     21404 => "00110101",
                     21405 => "10110101",
                     21406 => "01011000",
                     21407 => "01001001",
                     21408 => "11111111",
                     21409 => "00011000",
                     21410 => "01101001",
                     21411 => "00000001",
                     21412 => "10010101",
                     21413 => "01011000",
                     21414 => "11110110",
                     21415 => "10100000",
                     21416 => "10111101",
                     21417 => "00110100",
                     21418 => "00000100",
                     21419 => "10110100",
                     21420 => "01011000",
                     21421 => "00010000",
                     21422 => "00000011",
                     21423 => "10111101",
                     21424 => "00010111",
                     21425 => "00000100",
                     21426 => "10000101",
                     21427 => "00000000",
                     21428 => "10100101",
                     21429 => "00001001",
                     21430 => "01001010",
                     21431 => "10010000",
                     21432 => "00011001",
                     21433 => "10101101",
                     21434 => "01000111",
                     21435 => "00000111",
                     21436 => "11010000",
                     21437 => "00010100",
                     21438 => "10110101",
                     21439 => "11001111",
                     21440 => "00011000",
                     21441 => "01110101",
                     21442 => "01011000",
                     21443 => "10010101",
                     21444 => "11001111",
                     21445 => "11000101",
                     21446 => "00000000",
                     21447 => "11010000",
                     21448 => "00001001",
                     21449 => "10101001",
                     21450 => "00000000",
                     21451 => "10010101",
                     21452 => "10100000",
                     21453 => "10101001",
                     21454 => "01000000",
                     21455 => "10011101",
                     21456 => "10001010",
                     21457 => "00000111",
                     21458 => "10101001",
                     21459 => "00100000",
                     21460 => "10011101",
                     21461 => "11000101",
                     21462 => "00000011",
                     21463 => "01100000",
                     21464 => "10000101",
                     21465 => "00000111",
                     21466 => "10110101",
                     21467 => "00110100",
                     21468 => "11010000",
                     21469 => "00001110",
                     21470 => "10100000",
                     21471 => "00011000",
                     21472 => "10110101",
                     21473 => "01011000",
                     21474 => "00011000",
                     21475 => "01100101",
                     21476 => "00000111",
                     21477 => "10010101",
                     21478 => "01011000",
                     21479 => "10110101",
                     21480 => "10100000",
                     21481 => "01101001",
                     21482 => "00000000",
                     21483 => "01100000",
                     21484 => "10100000",
                     21485 => "00001000",
                     21486 => "10110101",
                     21487 => "01011000",
                     21488 => "00111000",
                     21489 => "11100101",
                     21490 => "00000111",
                     21491 => "10010101",
                     21492 => "01011000",
                     21493 => "10110101",
                     21494 => "10100000",
                     21495 => "11101001",
                     21496 => "00000000",
                     21497 => "01100000",
                     21498 => "10110101",
                     21499 => "10110110",
                     21500 => "11001001",
                     21501 => "00000011",
                     21502 => "11010000",
                     21503 => "00000011",
                     21504 => "01001100",
                     21505 => "10011110",
                     21506 => "11001001",
                     21507 => "10110101",
                     21508 => "00011110",
                     21509 => "00010000",
                     21510 => "00000001",
                     21511 => "01100000",
                     21512 => "10101000",
                     21513 => "10111101",
                     21514 => "10100010",
                     21515 => "00000011",
                     21516 => "10000101",
                     21517 => "00000000",
                     21518 => "10110101",
                     21519 => "01000110",
                     21520 => "11110000",
                     21521 => "00000011",
                     21522 => "01001100",
                     21523 => "10000011",
                     21524 => "11010101",
                     21525 => "10101001",
                     21526 => "00101101",
                     21527 => "11010101",
                     21528 => "11001111",
                     21529 => "10010000",
                     21530 => "00001111",
                     21531 => "11000100",
                     21532 => "00000000",
                     21533 => "11110000",
                     21534 => "00001000",
                     21535 => "00011000",
                     21536 => "01101001",
                     21537 => "00000010",
                     21538 => "10010101",
                     21539 => "11001111",
                     21540 => "01001100",
                     21541 => "01111001",
                     21542 => "11010101",
                     21543 => "01001100",
                     21544 => "01100000",
                     21545 => "11010101",
                     21546 => "11011001",
                     21547 => "11001111",
                     21548 => "00000000",
                     21549 => "10010000",
                     21550 => "00001101",
                     21551 => "11100100",
                     21552 => "00000000",
                     21553 => "11110000",
                     21554 => "11110100",
                     21555 => "00011000",
                     21556 => "01101001",
                     21557 => "00000010",
                     21558 => "10011001",
                     21559 => "11001111",
                     21560 => "00000000",
                     21561 => "01001100",
                     21562 => "01111001",
                     21563 => "11010101",
                     21564 => "10110101",
                     21565 => "11001111",
                     21566 => "01001000",
                     21567 => "10111101",
                     21568 => "10100010",
                     21569 => "00000011",
                     21570 => "00010000",
                     21571 => "00011000",
                     21572 => "10111101",
                     21573 => "00110100",
                     21574 => "00000100",
                     21575 => "00011000",
                     21576 => "01101001",
                     21577 => "00000101",
                     21578 => "10000101",
                     21579 => "00000000",
                     21580 => "10110101",
                     21581 => "10100000",
                     21582 => "01101001",
                     21583 => "00000000",
                     21584 => "00110000",
                     21585 => "00011010",
                     21586 => "11010000",
                     21587 => "00001100",
                     21588 => "10100101",
                     21589 => "00000000",
                     21590 => "11001001",
                     21591 => "00001011",
                     21592 => "10010000",
                     21593 => "00001100",
                     21594 => "10110000",
                     21595 => "00000100",
                     21596 => "11000101",
                     21597 => "00001000",
                     21598 => "11110000",
                     21599 => "00001100",
                     21600 => "00100000",
                     21601 => "10111100",
                     21602 => "10111111",
                     21603 => "01001100",
                     21604 => "01101111",
                     21605 => "11010100",
                     21606 => "00100000",
                     21607 => "01111001",
                     21608 => "11010101",
                     21609 => "01001100",
                     21610 => "01101111",
                     21611 => "11010100",
                     21612 => "00100000",
                     21613 => "10111001",
                     21614 => "10111111",
                     21615 => "10110100",
                     21616 => "00011110",
                     21617 => "01101000",
                     21618 => "00111000",
                     21619 => "11110101",
                     21620 => "11001111",
                     21621 => "00011000",
                     21622 => "01111001",
                     21623 => "11001111",
                     21624 => "00000000",
                     21625 => "10011001",
                     21626 => "11001111",
                     21627 => "00000000",
                     21628 => "10111101",
                     21629 => "10100010",
                     21630 => "00000011",
                     21631 => "00110000",
                     21632 => "00000100",
                     21633 => "10101010",
                     21634 => "00100000",
                     21635 => "00100011",
                     21636 => "11011100",
                     21637 => "10100100",
                     21638 => "00001000",
                     21639 => "10111001",
                     21640 => "10100000",
                     21641 => "00000000",
                     21642 => "00011001",
                     21643 => "00110100",
                     21644 => "00000100",
                     21645 => "11110000",
                     21646 => "01110111",
                     21647 => "10101110",
                     21648 => "00000000",
                     21649 => "00000011",
                     21650 => "11100000",
                     21651 => "00100000",
                     21652 => "10110000",
                     21653 => "01110000",
                     21654 => "10111001",
                     21655 => "10100000",
                     21656 => "00000000",
                     21657 => "01001000",
                     21658 => "01001000",
                     21659 => "00100000",
                     21660 => "00001001",
                     21661 => "11010101",
                     21662 => "10100101",
                     21663 => "00000001",
                     21664 => "10011101",
                     21665 => "00000001",
                     21666 => "00000011",
                     21667 => "10100101",
                     21668 => "00000000",
                     21669 => "10011101",
                     21670 => "00000010",
                     21671 => "00000011",
                     21672 => "10101001",
                     21673 => "00000010",
                     21674 => "10011101",
                     21675 => "00000011",
                     21676 => "00000011",
                     21677 => "10111001",
                     21678 => "10100000",
                     21679 => "00000000",
                     21680 => "00110000",
                     21681 => "00001101",
                     21682 => "10101001",
                     21683 => "10100010",
                     21684 => "10011101",
                     21685 => "00000100",
                     21686 => "00000011",
                     21687 => "10101001",
                     21688 => "10100011",
                     21689 => "10011101",
                     21690 => "00000101",
                     21691 => "00000011",
                     21692 => "01001100",
                     21693 => "11000111",
                     21694 => "11010100",
                     21695 => "10101001",
                     21696 => "00100100",
                     21697 => "10011101",
                     21698 => "00000100",
                     21699 => "00000011",
                     21700 => "10011101",
                     21701 => "00000101",
                     21702 => "00000011",
                     21703 => "10111001",
                     21704 => "00011110",
                     21705 => "00000000",
                     21706 => "10101000",
                     21707 => "01101000",
                     21708 => "01001001",
                     21709 => "11111111",
                     21710 => "00100000",
                     21711 => "00001001",
                     21712 => "11010101",
                     21713 => "10100101",
                     21714 => "00000001",
                     21715 => "10011101",
                     21716 => "00000110",
                     21717 => "00000011",
                     21718 => "10100101",
                     21719 => "00000000",
                     21720 => "10011101",
                     21721 => "00000111",
                     21722 => "00000011",
                     21723 => "10101001",
                     21724 => "00000010",
                     21725 => "10011101",
                     21726 => "00001000",
                     21727 => "00000011",
                     21728 => "01101000",
                     21729 => "00010000",
                     21730 => "00001101",
                     21731 => "10101001",
                     21732 => "10100010",
                     21733 => "10011101",
                     21734 => "00001001",
                     21735 => "00000011",
                     21736 => "10101001",
                     21737 => "10100011",
                     21738 => "10011101",
                     21739 => "00001010",
                     21740 => "00000011",
                     21741 => "01001100",
                     21742 => "11111000",
                     21743 => "11010100",
                     21744 => "10101001",
                     21745 => "00100100",
                     21746 => "10011101",
                     21747 => "00001001",
                     21748 => "00000011",
                     21749 => "10011101",
                     21750 => "00001010",
                     21751 => "00000011",
                     21752 => "10101001",
                     21753 => "00000000",
                     21754 => "10011101",
                     21755 => "00001011",
                     21756 => "00000011",
                     21757 => "10101101",
                     21758 => "00000000",
                     21759 => "00000011",
                     21760 => "00011000",
                     21761 => "01101001",
                     21762 => "00001010",
                     21763 => "10001101",
                     21764 => "00000000",
                     21765 => "00000011",
                     21766 => "10100110",
                     21767 => "00001000",
                     21768 => "01100000",
                     21769 => "01001000",
                     21770 => "10111001",
                     21771 => "10000111",
                     21772 => "00000000",
                     21773 => "00011000",
                     21774 => "01101001",
                     21775 => "00001000",
                     21776 => "10101110",
                     21777 => "11001100",
                     21778 => "00000110",
                     21779 => "11010000",
                     21780 => "00000011",
                     21781 => "00011000",
                     21782 => "01101001",
                     21783 => "00010000",
                     21784 => "01001000",
                     21785 => "10111001",
                     21786 => "01101110",
                     21787 => "00000000",
                     21788 => "01101001",
                     21789 => "00000000",
                     21790 => "10000101",
                     21791 => "00000010",
                     21792 => "01101000",
                     21793 => "00101001",
                     21794 => "11110000",
                     21795 => "01001010",
                     21796 => "01001010",
                     21797 => "01001010",
                     21798 => "10000101",
                     21799 => "00000000",
                     21800 => "10110110",
                     21801 => "11001111",
                     21802 => "01101000",
                     21803 => "00010000",
                     21804 => "00000101",
                     21805 => "10001010",
                     21806 => "00011000",
                     21807 => "01101001",
                     21808 => "00001000",
                     21809 => "10101010",
                     21810 => "10001010",
                     21811 => "10101110",
                     21812 => "00000000",
                     21813 => "00000011",
                     21814 => "00001010",
                     21815 => "00101010",
                     21816 => "01001000",
                     21817 => "00101010",
                     21818 => "00101001",
                     21819 => "00000011",
                     21820 => "00001001",
                     21821 => "00100000",
                     21822 => "10000101",
                     21823 => "00000001",
                     21824 => "10100101",
                     21825 => "00000010",
                     21826 => "00101001",
                     21827 => "00000001",
                     21828 => "00001010",
                     21829 => "00001010",
                     21830 => "00000101",
                     21831 => "00000001",
                     21832 => "10000101",
                     21833 => "00000001",
                     21834 => "01101000",
                     21835 => "00101001",
                     21836 => "11100000",
                     21837 => "00011000",
                     21838 => "01100101",
                     21839 => "00000000",
                     21840 => "10000101",
                     21841 => "00000000",
                     21842 => "10111001",
                     21843 => "11001111",
                     21844 => "00000000",
                     21845 => "11001001",
                     21846 => "11101000",
                     21847 => "10010000",
                     21848 => "00000110",
                     21849 => "10100101",
                     21850 => "00000000",
                     21851 => "00101001",
                     21852 => "10111111",
                     21853 => "10000101",
                     21854 => "00000000",
                     21855 => "01100000",
                     21856 => "10011000",
                     21857 => "10101010",
                     21858 => "00100000",
                     21859 => "10110110",
                     21860 => "11110001",
                     21861 => "10101001",
                     21862 => "00000110",
                     21863 => "00100000",
                     21864 => "00010011",
                     21865 => "11011010",
                     21866 => "10101101",
                     21867 => "10101101",
                     21868 => "00000011",
                     21869 => "10011101",
                     21870 => "00010111",
                     21871 => "00000001",
                     21872 => "10100101",
                     21873 => "11001110",
                     21874 => "10011101",
                     21875 => "00011110",
                     21876 => "00000001",
                     21877 => "10101001",
                     21878 => "00000001",
                     21879 => "10010101",
                     21880 => "01000110",
                     21881 => "00100000",
                     21882 => "01101001",
                     21883 => "11000011",
                     21884 => "10011001",
                     21885 => "10100000",
                     21886 => "00000000",
                     21887 => "10011001",
                     21888 => "00110100",
                     21889 => "00000100",
                     21890 => "01100000",
                     21891 => "10011000",
                     21892 => "01001000",
                     21893 => "00100000",
                     21894 => "01110000",
                     21895 => "10111111",
                     21896 => "01101000",
                     21897 => "10101010",
                     21898 => "00100000",
                     21899 => "01110000",
                     21900 => "10111111",
                     21901 => "10100110",
                     21902 => "00001000",
                     21903 => "10111101",
                     21904 => "10100010",
                     21905 => "00000011",
                     21906 => "00110000",
                     21907 => "00000100",
                     21908 => "10101010",
                     21909 => "00100000",
                     21910 => "00100011",
                     21911 => "11011100",
                     21912 => "10100110",
                     21913 => "00001000",
                     21914 => "01100000",
                     21915 => "10110101",
                     21916 => "10100000",
                     21917 => "00011101",
                     21918 => "00110100",
                     21919 => "00000100",
                     21920 => "11010000",
                     21921 => "00010101",
                     21922 => "10011101",
                     21923 => "00010111",
                     21924 => "00000100",
                     21925 => "10110101",
                     21926 => "11001111",
                     21927 => "11011101",
                     21928 => "00000001",
                     21929 => "00000100",
                     21930 => "10110000",
                     21931 => "00001011",
                     21932 => "10100101",
                     21933 => "00001001",
                     21934 => "00101001",
                     21935 => "00000111",
                     21936 => "11010000",
                     21937 => "00000010",
                     21938 => "11110110",
                     21939 => "11001111",
                     21940 => "01001100",
                     21941 => "11000110",
                     21942 => "11010101",
                     21943 => "10110101",
                     21944 => "11001111",
                     21945 => "11010101",
                     21946 => "01011000",
                     21947 => "10010000",
                     21948 => "00000110",
                     21949 => "00100000",
                     21950 => "10111100",
                     21951 => "10111111",
                     21952 => "01001100",
                     21953 => "11000110",
                     21954 => "11010101",
                     21955 => "00100000",
                     21956 => "10111001",
                     21957 => "10111111",
                     21958 => "10111101",
                     21959 => "10100010",
                     21960 => "00000011",
                     21961 => "00110000",
                     21962 => "00000011",
                     21963 => "00100000",
                     21964 => "00100011",
                     21965 => "11011100",
                     21966 => "01100000",
                     21967 => "10101001",
                     21968 => "00001110",
                     21969 => "00100000",
                     21970 => "01001101",
                     21971 => "11001011",
                     21972 => "00100000",
                     21973 => "01101100",
                     21974 => "11001011",
                     21975 => "10111101",
                     21976 => "10100010",
                     21977 => "00000011",
                     21978 => "00110000",
                     21979 => "00011100",
                     21980 => "10100101",
                     21981 => "10000110",
                     21982 => "00011000",
                     21983 => "01100101",
                     21984 => "00000000",
                     21985 => "10000101",
                     21986 => "10000110",
                     21987 => "10100101",
                     21988 => "01101101",
                     21989 => "10100100",
                     21990 => "00000000",
                     21991 => "00110000",
                     21992 => "00000101",
                     21993 => "01101001",
                     21994 => "00000000",
                     21995 => "01001100",
                     21996 => "11110000",
                     21997 => "11010101",
                     21998 => "11101001",
                     21999 => "00000000",
                     22000 => "10000101",
                     22001 => "01101101",
                     22002 => "10001100",
                     22003 => "10100001",
                     22004 => "00000011",
                     22005 => "00100000",
                     22006 => "00100011",
                     22007 => "11011100",
                     22008 => "01100000",
                     22009 => "10111101",
                     22010 => "10100010",
                     22011 => "00000011",
                     22012 => "00110000",
                     22013 => "00000110",
                     22014 => "00100000",
                     22015 => "10001101",
                     22016 => "10111111",
                     22017 => "00100000",
                     22018 => "00100011",
                     22019 => "11011100",
                     22020 => "01100000",
                     22021 => "00100000",
                     22022 => "00000111",
                     22023 => "10111111",
                     22024 => "10000101",
                     22025 => "00000000",
                     22026 => "10111101",
                     22027 => "10100010",
                     22028 => "00000011",
                     22029 => "00110000",
                     22030 => "00000111",
                     22031 => "10101001",
                     22032 => "00010011",
                     22033 => "10010101",
                     22034 => "01011000",
                     22035 => "00100000",
                     22036 => "11011100",
                     22037 => "11010101",
                     22038 => "01100000",
                     22039 => "00100000",
                     22040 => "00100011",
                     22041 => "11010110",
                     22042 => "01001100",
                     22043 => "11000110",
                     22044 => "11010101",
                     22045 => "00100000",
                     22046 => "00100011",
                     22047 => "11010110",
                     22048 => "01001100",
                     22049 => "00111001",
                     22050 => "11010110",
                     22051 => "10101101",
                     22052 => "01000111",
                     22053 => "00000111",
                     22054 => "11010000",
                     22055 => "00011001",
                     22056 => "10111101",
                     22057 => "00010111",
                     22058 => "00000100",
                     22059 => "00011000",
                     22060 => "01111101",
                     22061 => "00110100",
                     22062 => "00000100",
                     22063 => "10011101",
                     22064 => "00010111",
                     22065 => "00000100",
                     22066 => "10110101",
                     22067 => "11001111",
                     22068 => "01110101",
                     22069 => "10100000",
                     22070 => "10010101",
                     22071 => "11001111",
                     22072 => "01100000",
                     22073 => "10111101",
                     22074 => "10100010",
                     22075 => "00000011",
                     22076 => "11110000",
                     22077 => "00000011",
                     22078 => "00100000",
                     22079 => "00011011",
                     22080 => "11011100",
                     22081 => "01100000",
                     22082 => "10110101",
                     22083 => "00010110",
                     22084 => "11001001",
                     22085 => "00010100",
                     22086 => "11110000",
                     22087 => "01010101",
                     22088 => "10101101",
                     22089 => "00011100",
                     22090 => "00000111",
                     22091 => "10110100",
                     22092 => "00010110",
                     22093 => "11000000",
                     22094 => "00000101",
                     22095 => "11110000",
                     22096 => "00000100",
                     22097 => "11000000",
                     22098 => "00001101",
                     22099 => "11010000",
                     22100 => "00000010",
                     22101 => "01101001",
                     22102 => "00111000",
                     22103 => "11101001",
                     22104 => "01001000",
                     22105 => "10000101",
                     22106 => "00000001",
                     22107 => "10101101",
                     22108 => "00011010",
                     22109 => "00000111",
                     22110 => "11101001",
                     22111 => "00000000",
                     22112 => "10000101",
                     22113 => "00000000",
                     22114 => "10101101",
                     22115 => "00011101",
                     22116 => "00000111",
                     22117 => "01101001",
                     22118 => "01001000",
                     22119 => "10000101",
                     22120 => "00000011",
                     22121 => "10101101",
                     22122 => "00011011",
                     22123 => "00000111",
                     22124 => "01101001",
                     22125 => "00000000",
                     22126 => "10000101",
                     22127 => "00000010",
                     22128 => "10110101",
                     22129 => "10000111",
                     22130 => "11000101",
                     22131 => "00000001",
                     22132 => "10110101",
                     22133 => "01101110",
                     22134 => "11100101",
                     22135 => "00000000",
                     22136 => "00110000",
                     22137 => "00100000",
                     22138 => "10110101",
                     22139 => "10000111",
                     22140 => "11000101",
                     22141 => "00000011",
                     22142 => "10110101",
                     22143 => "01101110",
                     22144 => "11100101",
                     22145 => "00000010",
                     22146 => "00110000",
                     22147 => "00011001",
                     22148 => "10110101",
                     22149 => "00011110",
                     22150 => "11001001",
                     22151 => "00000101",
                     22152 => "11110000",
                     22153 => "00010011",
                     22154 => "11000000",
                     22155 => "00001101",
                     22156 => "11110000",
                     22157 => "00001111",
                     22158 => "11000000",
                     22159 => "00110000",
                     22160 => "11110000",
                     22161 => "00001011",
                     22162 => "11000000",
                     22163 => "00110001",
                     22164 => "11110000",
                     22165 => "00000111",
                     22166 => "11000000",
                     22167 => "00110010",
                     22168 => "11110000",
                     22169 => "00000011",
                     22170 => "00100000",
                     22171 => "10011110",
                     22172 => "11001001",
                     22173 => "01100000",
                     22174 => "11111111",
                     22175 => "11111111",
                     22176 => "11111111",
                     22177 => "11111111",
                     22178 => "11111111",
                     22179 => "11111111",
                     22180 => "11111111",
                     22181 => "11111111",
                     22182 => "11111111",
                     22183 => "11111111",
                     22184 => "11111111",
                     22185 => "11111111",
                     22186 => "11111111",
                     22187 => "11111111",
                     22188 => "11111111",
                     22189 => "11111111",
                     22190 => "11111111",
                     22191 => "11111111",
                     22192 => "11111111",
                     22193 => "11111111",
                     22194 => "11111111",
                     22195 => "11111111",
                     22196 => "11111111",
                     22197 => "11111111",
                     22198 => "11111111",
                     22199 => "11111111",
                     22200 => "11111111",
                     22201 => "11111111",
                     22202 => "11111111",
                     22203 => "11111111",
                     22204 => "11111111",
                     22205 => "11111111",
                     22206 => "11111111",
                     22207 => "11111111",
                     22208 => "11111111",
                     22209 => "11111111",
                     22210 => "11111111",
                     22211 => "11111111",
                     22212 => "11111111",
                     22213 => "11111111",
                     22214 => "11111111",
                     22215 => "11111111",
                     22216 => "11111111",
                     22217 => "11111111",
                     22218 => "11111111",
                     22219 => "11111111",
                     22220 => "11111111",
                     22221 => "11111111",
                     22222 => "11111111",
                     22223 => "11111111",
                     22224 => "11111111",
                     22225 => "11111111",
                     22226 => "11111111",
                     22227 => "11111111",
                     22228 => "11111111",
                     22229 => "11111111",
                     22230 => "11111111",
                     22231 => "11111111",
                     22232 => "11111111",
                     22233 => "10110101",
                     22234 => "00100100",
                     22235 => "11110000",
                     22236 => "01010110",
                     22237 => "00001010",
                     22238 => "10110000",
                     22239 => "01010011",
                     22240 => "10100101",
                     22241 => "00001001",
                     22242 => "01001010",
                     22243 => "10110000",
                     22244 => "01001110",
                     22245 => "10001010",
                     22246 => "00001010",
                     22247 => "00001010",
                     22248 => "00011000",
                     22249 => "01101001",
                     22250 => "00011100",
                     22251 => "10101000",
                     22252 => "10100010",
                     22253 => "00000100",
                     22254 => "10000110",
                     22255 => "00000001",
                     22256 => "10011000",
                     22257 => "01001000",
                     22258 => "10110101",
                     22259 => "00011110",
                     22260 => "00101001",
                     22261 => "00100000",
                     22262 => "11010000",
                     22263 => "00110100",
                     22264 => "10110101",
                     22265 => "00001111",
                     22266 => "11110000",
                     22267 => "00110000",
                     22268 => "10110101",
                     22269 => "00010110",
                     22270 => "11001001",
                     22271 => "00100100",
                     22272 => "10010000",
                     22273 => "00000100",
                     22274 => "11001001",
                     22275 => "00101011",
                     22276 => "10010000",
                     22277 => "00100110",
                     22278 => "11001001",
                     22279 => "00000110",
                     22280 => "11010000",
                     22281 => "00000110",
                     22282 => "10110101",
                     22283 => "00011110",
                     22284 => "11001001",
                     22285 => "00000010",
                     22286 => "10110000",
                     22287 => "00011100",
                     22288 => "10111101",
                     22289 => "11011000",
                     22290 => "00000011",
                     22291 => "11010000",
                     22292 => "00010111",
                     22293 => "10001010",
                     22294 => "00001010",
                     22295 => "00001010",
                     22296 => "00011000",
                     22297 => "01101001",
                     22298 => "00000100",
                     22299 => "10101010",
                     22300 => "00100000",
                     22301 => "00101111",
                     22302 => "11100011",
                     22303 => "10100110",
                     22304 => "00001000",
                     22305 => "10010000",
                     22306 => "00001001",
                     22307 => "10101001",
                     22308 => "10000000",
                     22309 => "10010101",
                     22310 => "00100100",
                     22311 => "10100110",
                     22312 => "00000001",
                     22313 => "00100000",
                     22314 => "00111110",
                     22315 => "11010111",
                     22316 => "01101000",
                     22317 => "10101000",
                     22318 => "10100110",
                     22319 => "00000001",
                     22320 => "11001010",
                     22321 => "00010000",
                     22322 => "10111011",
                     22323 => "10100110",
                     22324 => "00001000",
                     22325 => "01100000",
                     22326 => "00000110",
                     22327 => "00000000",
                     22328 => "00000010",
                     22329 => "00010010",
                     22330 => "00010001",
                     22331 => "00000111",
                     22332 => "00000101",
                     22333 => "00101101",
                     22334 => "00100000",
                     22335 => "01011001",
                     22336 => "11110001",
                     22337 => "10100110",
                     22338 => "00000001",
                     22339 => "10110101",
                     22340 => "00001111",
                     22341 => "00010000",
                     22342 => "00001011",
                     22343 => "00101001",
                     22344 => "00001111",
                     22345 => "10101010",
                     22346 => "10110101",
                     22347 => "00010110",
                     22348 => "11001001",
                     22349 => "00101101",
                     22350 => "11110000",
                     22351 => "00001100",
                     22352 => "10100110",
                     22353 => "00000001",
                     22354 => "10110101",
                     22355 => "00010110",
                     22356 => "11001001",
                     22357 => "00000010",
                     22358 => "11110000",
                     22359 => "01101011",
                     22360 => "11001001",
                     22361 => "00101101",
                     22362 => "11010000",
                     22363 => "00101101",
                     22364 => "11001110",
                     22365 => "10000011",
                     22366 => "00000100",
                     22367 => "11010000",
                     22368 => "01100010",
                     22369 => "00100000",
                     22370 => "01101001",
                     22371 => "11000011",
                     22372 => "10010101",
                     22373 => "01011000",
                     22374 => "10001101",
                     22375 => "11001011",
                     22376 => "00000110",
                     22377 => "10101001",
                     22378 => "11111110",
                     22379 => "10010101",
                     22380 => "10100000",
                     22381 => "10101100",
                     22382 => "01011111",
                     22383 => "00000111",
                     22384 => "10111001",
                     22385 => "00110110",
                     22386 => "11010111",
                     22387 => "10010101",
                     22388 => "00010110",
                     22389 => "10101001",
                     22390 => "00100000",
                     22391 => "11000000",
                     22392 => "00000011",
                     22393 => "10110000",
                     22394 => "00000010",
                     22395 => "00001001",
                     22396 => "00000011",
                     22397 => "10010101",
                     22398 => "00011110",
                     22399 => "10101001",
                     22400 => "10000000",
                     22401 => "10000101",
                     22402 => "11111110",
                     22403 => "10100110",
                     22404 => "00000001",
                     22405 => "10101001",
                     22406 => "00001001",
                     22407 => "11010000",
                     22408 => "00110011",
                     22409 => "11001001",
                     22410 => "00001000",
                     22411 => "11110000",
                     22412 => "00110110",
                     22413 => "11001001",
                     22414 => "00001100",
                     22415 => "11110000",
                     22416 => "00110010",
                     22417 => "11001001",
                     22418 => "00010101",
                     22419 => "10110000",
                     22420 => "00101110",
                     22421 => "10110101",
                     22422 => "00010110",
                     22423 => "11001001",
                     22424 => "00001101",
                     22425 => "11010000",
                     22426 => "00000110",
                     22427 => "10110101",
                     22428 => "11001111",
                     22429 => "01101001",
                     22430 => "00011000",
                     22431 => "10010101",
                     22432 => "11001111",
                     22433 => "00100000",
                     22434 => "00100011",
                     22435 => "11100000",
                     22436 => "10110101",
                     22437 => "00011110",
                     22438 => "00101001",
                     22439 => "00011111",
                     22440 => "00001001",
                     22441 => "00100000",
                     22442 => "10010101",
                     22443 => "00011110",
                     22444 => "10101001",
                     22445 => "00000010",
                     22446 => "10110100",
                     22447 => "00010110",
                     22448 => "11000000",
                     22449 => "00000101",
                     22450 => "11010000",
                     22451 => "00000010",
                     22452 => "10101001",
                     22453 => "00000110",
                     22454 => "11000000",
                     22455 => "00000110",
                     22456 => "11010000",
                     22457 => "00000010",
                     22458 => "10101001",
                     22459 => "00000001",
                     22460 => "00100000",
                     22461 => "00010011",
                     22462 => "11011010",
                     22463 => "10101001",
                     22464 => "00001000",
                     22465 => "10000101",
                     22466 => "11111111",
                     22467 => "01100000",
                     22468 => "10100101",
                     22469 => "00001001",
                     22470 => "01001010",
                     22471 => "10010000",
                     22472 => "00110110",
                     22473 => "10101101",
                     22474 => "01000111",
                     22475 => "00000111",
                     22476 => "00001101",
                     22477 => "11010110",
                     22478 => "00000011",
                     22479 => "11010000",
                     22480 => "00101110",
                     22481 => "10001010",
                     22482 => "00001010",
                     22483 => "00001010",
                     22484 => "00011000",
                     22485 => "01101001",
                     22486 => "00100100",
                     22487 => "10101000",
                     22488 => "00100000",
                     22489 => "00101101",
                     22490 => "11100011",
                     22491 => "10100110",
                     22492 => "00001000",
                     22493 => "10010000",
                     22494 => "00011011",
                     22495 => "10111101",
                     22496 => "10111110",
                     22497 => "00000110",
                     22498 => "11010000",
                     22499 => "00011011",
                     22500 => "10101001",
                     22501 => "00000001",
                     22502 => "10011101",
                     22503 => "10111110",
                     22504 => "00000110",
                     22505 => "10110101",
                     22506 => "01100100",
                     22507 => "01001001",
                     22508 => "11111111",
                     22509 => "00011000",
                     22510 => "01101001",
                     22511 => "00000001",
                     22512 => "10010101",
                     22513 => "01100100",
                     22514 => "10101101",
                     22515 => "10011111",
                     22516 => "00000111",
                     22517 => "11010000",
                     22518 => "00001000",
                     22519 => "01001100",
                     22520 => "00101101",
                     22521 => "11011001",
                     22522 => "10101001",
                     22523 => "00000000",
                     22524 => "10011101",
                     22525 => "10111110",
                     22526 => "00000110",
                     22527 => "01100000",
                     22528 => "00100000",
                     22529 => "10011110",
                     22530 => "11001001",
                     22531 => "10101001",
                     22532 => "00000110",
                     22533 => "00100000",
                     22534 => "00010011",
                     22535 => "11011010",
                     22536 => "10101001",
                     22537 => "00100000",
                     22538 => "10000101",
                     22539 => "11111110",
                     22540 => "10100101",
                     22541 => "00111001",
                     22542 => "11001001",
                     22543 => "00000010",
                     22544 => "10010000",
                     22545 => "00001110",
                     22546 => "11001001",
                     22547 => "00000011",
                     22548 => "11110000",
                     22549 => "00100100",
                     22550 => "10101001",
                     22551 => "00100011",
                     22552 => "10001101",
                     22553 => "10011111",
                     22554 => "00000111",
                     22555 => "10101001",
                     22556 => "01000000",
                     22557 => "10000101",
                     22558 => "11111011",
                     22559 => "01100000",
                     22560 => "10101101",
                     22561 => "01010110",
                     22562 => "00000111",
                     22563 => "11110000",
                     22564 => "00011011",
                     22565 => "11001001",
                     22566 => "00000001",
                     22567 => "11010000",
                     22568 => "00100011",
                     22569 => "10100110",
                     22570 => "00001000",
                     22571 => "10101001",
                     22572 => "00000010",
                     22573 => "10001101",
                     22574 => "01010110",
                     22575 => "00000111",
                     22576 => "00100000",
                     22577 => "11110001",
                     22578 => "10000101",
                     22579 => "10100110",
                     22580 => "00001000",
                     22581 => "10101001",
                     22582 => "00001100",
                     22583 => "01001100",
                     22584 => "01000111",
                     22585 => "11011000",
                     22586 => "10101001",
                     22587 => "00001011",
                     22588 => "10011101",
                     22589 => "00010000",
                     22590 => "00000001",
                     22591 => "01100000",
                     22592 => "10101001",
                     22593 => "00000001",
                     22594 => "10001101",
                     22595 => "01010110",
                     22596 => "00000111",
                     22597 => "10101001",
                     22598 => "00001001",
                     22599 => "10100000",
                     22600 => "00000000",
                     22601 => "00100000",
                     22602 => "01001010",
                     22603 => "11011001",
                     22604 => "01100000",
                     22605 => "00011000",
                     22606 => "11101000",
                     22607 => "00111000",
                     22608 => "11001000",
                     22609 => "00001000",
                     22610 => "11111000",
                     22611 => "10100101",
                     22612 => "00001001",
                     22613 => "01001010",
                     22614 => "10110000",
                     22615 => "11110100",
                     22616 => "00100000",
                     22617 => "01000011",
                     22618 => "11011100",
                     22619 => "10110000",
                     22620 => "00100011",
                     22621 => "10111101",
                     22622 => "11011000",
                     22623 => "00000011",
                     22624 => "11010000",
                     22625 => "00011110",
                     22626 => "10100101",
                     22627 => "00001110",
                     22628 => "11001001",
                     22629 => "00001000",
                     22630 => "11010000",
                     22631 => "00011000",
                     22632 => "10110101",
                     22633 => "00011110",
                     22634 => "00101001",
                     22635 => "00100000",
                     22636 => "11010000",
                     22637 => "00010010",
                     22638 => "00100000",
                     22639 => "01010100",
                     22640 => "11011100",
                     22641 => "00100000",
                     22642 => "00101101",
                     22643 => "11100011",
                     22644 => "10100110",
                     22645 => "00001000",
                     22646 => "10110000",
                     22647 => "00001001",
                     22648 => "10111101",
                     22649 => "10010001",
                     22650 => "00000100",
                     22651 => "00101001",
                     22652 => "11111110",
                     22653 => "10011101",
                     22654 => "10010001",
                     22655 => "00000100",
                     22656 => "01100000",
                     22657 => "10110100",
                     22658 => "00010110",
                     22659 => "11000000",
                     22660 => "00101110",
                     22661 => "11010000",
                     22662 => "00000011",
                     22663 => "01001100",
                     22664 => "00000000",
                     22665 => "11011000",
                     22666 => "10101101",
                     22667 => "10011111",
                     22668 => "00000111",
                     22669 => "11110000",
                     22670 => "00000110",
                     22671 => "01001100",
                     22672 => "10010101",
                     22673 => "11010111",
                     22674 => "00001010",
                     22675 => "00000110",
                     22676 => "00000100",
                     22677 => "10111101",
                     22678 => "10010001",
                     22679 => "00000100",
                     22680 => "00101001",
                     22681 => "00000001",
                     22682 => "00011101",
                     22683 => "11011000",
                     22684 => "00000011",
                     22685 => "11010000",
                     22686 => "01011001",
                     22687 => "10101001",
                     22688 => "00000001",
                     22689 => "00011101",
                     22690 => "10010001",
                     22691 => "00000100",
                     22692 => "10011101",
                     22693 => "10010001",
                     22694 => "00000100",
                     22695 => "11000000",
                     22696 => "00010010",
                     22697 => "11110000",
                     22698 => "01001110",
                     22699 => "11000000",
                     22700 => "00001101",
                     22701 => "11110000",
                     22702 => "01111110",
                     22703 => "11000000",
                     22704 => "00001100",
                     22705 => "11110000",
                     22706 => "01111010",
                     22707 => "11000000",
                     22708 => "00110011",
                     22709 => "11110000",
                     22710 => "01000010",
                     22711 => "11000000",
                     22712 => "00010101",
                     22713 => "10110000",
                     22714 => "01110010",
                     22715 => "10101101",
                     22716 => "01001110",
                     22717 => "00000111",
                     22718 => "11110000",
                     22719 => "01101101",
                     22720 => "10110101",
                     22721 => "00011110",
                     22722 => "00001010",
                     22723 => "10110000",
                     22724 => "00110100",
                     22725 => "10110101",
                     22726 => "00011110",
                     22727 => "00101001",
                     22728 => "00000111",
                     22729 => "11001001",
                     22730 => "00000010",
                     22731 => "10010000",
                     22732 => "00101100",
                     22733 => "10110101",
                     22734 => "00010110",
                     22735 => "11001001",
                     22736 => "00000110",
                     22737 => "11110000",
                     22738 => "00100101",
                     22739 => "10101001",
                     22740 => "00001000",
                     22741 => "10000101",
                     22742 => "11111111",
                     22743 => "10110101",
                     22744 => "00011110",
                     22745 => "00001001",
                     22746 => "10000000",
                     22747 => "10010101",
                     22748 => "00011110",
                     22749 => "00100000",
                     22750 => "00000111",
                     22751 => "11011010",
                     22752 => "10111001",
                     22753 => "01001111",
                     22754 => "11011000",
                     22755 => "10010101",
                     22756 => "01011000",
                     22757 => "10101001",
                     22758 => "00000011",
                     22759 => "00011000",
                     22760 => "01101101",
                     22761 => "10000100",
                     22762 => "00000100",
                     22763 => "10111100",
                     22764 => "10010110",
                     22765 => "00000111",
                     22766 => "11000000",
                     22767 => "00000011",
                     22768 => "10110000",
                     22769 => "00000011",
                     22770 => "10111001",
                     22771 => "10010010",
                     22772 => "11011000",
                     22773 => "00100000",
                     22774 => "00010011",
                     22775 => "11011010",
                     22776 => "01100000",
                     22777 => "10100101",
                     22778 => "10011111",
                     22779 => "00110000",
                     22780 => "00000010",
                     22781 => "11010000",
                     22782 => "01101100",
                     22783 => "10101001",
                     22784 => "00010100",
                     22785 => "10110100",
                     22786 => "00010110",
                     22787 => "11000000",
                     22788 => "00010100",
                     22789 => "11010000",
                     22790 => "00000010",
                     22791 => "10101001",
                     22792 => "00000111",
                     22793 => "01100101",
                     22794 => "11001110",
                     22795 => "11010101",
                     22796 => "11001111",
                     22797 => "10010000",
                     22798 => "01011100",
                     22799 => "10101101",
                     22800 => "10010001",
                     22801 => "00000111",
                     22802 => "11010000",
                     22803 => "01010111",
                     22804 => "10101101",
                     22805 => "10011110",
                     22806 => "00000111",
                     22807 => "11010000",
                     22808 => "00111110",
                     22809 => "10101101",
                     22810 => "10101101",
                     22811 => "00000011",
                     22812 => "11001101",
                     22813 => "10101110",
                     22814 => "00000011",
                     22815 => "10010000",
                     22816 => "00000011",
                     22817 => "01001100",
                     22818 => "11111000",
                     22819 => "11011001",
                     22820 => "10110101",
                     22821 => "01000110",
                     22822 => "11001001",
                     22823 => "00000001",
                     22824 => "11010000",
                     22825 => "00000011",
                     22826 => "01001100",
                     22827 => "00000001",
                     22828 => "11011010",
                     22829 => "10101101",
                     22830 => "10011110",
                     22831 => "00000111",
                     22832 => "11010000",
                     22833 => "00100101",
                     22834 => "10101110",
                     22835 => "01010110",
                     22836 => "00000111",
                     22837 => "11110000",
                     22838 => "00100011",
                     22839 => "10001101",
                     22840 => "01010110",
                     22841 => "00000111",
                     22842 => "10101001",
                     22843 => "00001000",
                     22844 => "10001101",
                     22845 => "10011110",
                     22846 => "00000111",
                     22847 => "10101001",
                     22848 => "00010000",
                     22849 => "10000101",
                     22850 => "11111111",
                     22851 => "00100000",
                     22852 => "11110001",
                     22853 => "10000101",
                     22854 => "10101001",
                     22855 => "00001010",
                     22856 => "10100000",
                     22857 => "00000001",
                     22858 => "10000101",
                     22859 => "00001110",
                     22860 => "10000100",
                     22861 => "00011101",
                     22862 => "10100000",
                     22863 => "11111111",
                     22864 => "10001100",
                     22865 => "01000111",
                     22866 => "00000111",
                     22867 => "11001000",
                     22868 => "10001100",
                     22869 => "01110101",
                     22870 => "00000111",
                     22871 => "10100110",
                     22872 => "00001000",
                     22873 => "01100000",
                     22874 => "10000110",
                     22875 => "01010111",
                     22876 => "11101000",
                     22877 => "10000110",
                     22878 => "11111100",
                     22879 => "10101001",
                     22880 => "11111100",
                     22881 => "10000101",
                     22882 => "10011111",
                     22883 => "10101001",
                     22884 => "00001011",
                     22885 => "11010000",
                     22886 => "11100001",
                     22887 => "00000010",
                     22888 => "00000110",
                     22889 => "00000101",
                     22890 => "00000110",
                     22891 => "10110101",
                     22892 => "00010110",
                     22893 => "11001001",
                     22894 => "00010010",
                     22895 => "11110000",
                     22896 => "10111100",
                     22897 => "10101001",
                     22898 => "00000100",
                     22899 => "10000101",
                     22900 => "11111111",
                     22901 => "10110101",
                     22902 => "00010110",
                     22903 => "10100000",
                     22904 => "00000000",
                     22905 => "11001001",
                     22906 => "00010100",
                     22907 => "11110000",
                     22908 => "00011011",
                     22909 => "11001001",
                     22910 => "00001000",
                     22911 => "11110000",
                     22912 => "00010111",
                     22913 => "11001001",
                     22914 => "00110011",
                     22915 => "11110000",
                     22916 => "00010011",
                     22917 => "11001001",
                     22918 => "00001100",
                     22919 => "11110000",
                     22920 => "00001111",
                     22921 => "11001000",
                     22922 => "11001001",
                     22923 => "00000101",
                     22924 => "11110000",
                     22925 => "00001010",
                     22926 => "11001000",
                     22927 => "11001001",
                     22928 => "00010001",
                     22929 => "11110000",
                     22930 => "00000101",
                     22931 => "11001000",
                     22932 => "11001001",
                     22933 => "00000111",
                     22934 => "11010000",
                     22935 => "00011101",
                     22936 => "10111001",
                     22937 => "01100111",
                     22938 => "11011001",
                     22939 => "00100000",
                     22940 => "00010011",
                     22941 => "11011010",
                     22942 => "10110101",
                     22943 => "01000110",
                     22944 => "01001000",
                     22945 => "00100000",
                     22946 => "00110111",
                     22947 => "11100000",
                     22948 => "01101000",
                     22949 => "10010101",
                     22950 => "01000110",
                     22951 => "10101001",
                     22952 => "00100000",
                     22953 => "10010101",
                     22954 => "00011110",
                     22955 => "00100000",
                     22956 => "01101001",
                     22957 => "11000011",
                     22958 => "10010101",
                     22959 => "01011000",
                     22960 => "10101001",
                     22961 => "11111101",
                     22962 => "10000101",
                     22963 => "10011111",
                     22964 => "01100000",
                     22965 => "11001001",
                     22966 => "00001001",
                     22967 => "10010000",
                     22968 => "00011101",
                     22969 => "00101001",
                     22970 => "00000001",
                     22971 => "10010101",
                     22972 => "00010110",
                     22973 => "10100000",
                     22974 => "00000000",
                     22975 => "10010100",
                     22976 => "00011110",
                     22977 => "10101001",
                     22978 => "00000011",
                     22979 => "00100000",
                     22980 => "00010011",
                     22981 => "11011010",
                     22982 => "00100000",
                     22983 => "01101001",
                     22984 => "11000011",
                     22985 => "00100000",
                     22986 => "00000111",
                     22987 => "11011010",
                     22988 => "10111001",
                     22989 => "01010001",
                     22990 => "11011000",
                     22991 => "10010101",
                     22992 => "01011000",
                     22993 => "01001100",
                     22994 => "11110011",
                     22995 => "11011001",
                     22996 => "00001101",
                     22997 => "00001001",
                     22998 => "10101001",
                     22999 => "00000100",
                     23000 => "10010101",
                     23001 => "00011110",
                     23002 => "11101110",
                     23003 => "10000100",
                     23004 => "00000100",
                     23005 => "10101101",
                     23006 => "10000100",
                     23007 => "00000100",
                     23008 => "00011000",
                     23009 => "01101101",
                     23010 => "10010001",
                     23011 => "00000111",
                     23012 => "00100000",
                     23013 => "00010011",
                     23014 => "11011010",
                     23015 => "11101110",
                     23016 => "10010001",
                     23017 => "00000111",
                     23018 => "10101100",
                     23019 => "01101010",
                     23020 => "00000111",
                     23021 => "10111001",
                     23022 => "11010100",
                     23023 => "11011001",
                     23024 => "10011101",
                     23025 => "10010110",
                     23026 => "00000111",
                     23027 => "10101001",
                     23028 => "11111100",
                     23029 => "10000101",
                     23030 => "10011111",
                     23031 => "01100000",
                     23032 => "10110101",
                     23033 => "01000110",
                     23034 => "11001001",
                     23035 => "00000001",
                     23036 => "11010000",
                     23037 => "00000011",
                     23038 => "01001100",
                     23039 => "00101101",
                     23040 => "11011001",
                     23041 => "00100000",
                     23042 => "00011110",
                     23043 => "11011011",
                     23044 => "01001100",
                     23045 => "00101101",
                     23046 => "11011001",
                     23047 => "10100000",
                     23048 => "00000001",
                     23049 => "00100000",
                     23050 => "01001011",
                     23051 => "11100001",
                     23052 => "00010000",
                     23053 => "00000001",
                     23054 => "11001000",
                     23055 => "10010100",
                     23056 => "01000110",
                     23057 => "10001000",
                     23058 => "01100000",
                     23059 => "10011101",
                     23060 => "00010000",
                     23061 => "00000001",
                     23062 => "10101001",
                     23063 => "00110000",
                     23064 => "10011101",
                     23065 => "00101100",
                     23066 => "00000001",
                     23067 => "10110101",
                     23068 => "11001111",
                     23069 => "10011101",
                     23070 => "00011110",
                     23071 => "00000001",
                     23072 => "10101101",
                     23073 => "10101110",
                     23074 => "00000011",
                     23075 => "10011101",
                     23076 => "00010111",
                     23077 => "00000001",
                     23078 => "01100000",
                     23079 => "10000000",
                     23080 => "01000000",
                     23081 => "00100000",
                     23082 => "00010000",
                     23083 => "00001000",
                     23084 => "00000100",
                     23085 => "00000010",
                     23086 => "01111111",
                     23087 => "10111111",
                     23088 => "11011111",
                     23089 => "11101111",
                     23090 => "11110111",
                     23091 => "11111011",
                     23092 => "11111101",
                     23093 => "10100101",
                     23094 => "00001001",
                     23095 => "01001010",
                     23096 => "10010000",
                     23097 => "11101100",
                     23098 => "10101101",
                     23099 => "01001110",
                     23100 => "00000111",
                     23101 => "11110000",
                     23102 => "11100111",
                     23103 => "10110101",
                     23104 => "00010110",
                     23105 => "11001001",
                     23106 => "00010101",
                     23107 => "10110000",
                     23108 => "01101110",
                     23109 => "11001001",
                     23110 => "00010001",
                     23111 => "11110000",
                     23112 => "01101010",
                     23113 => "11001001",
                     23114 => "00001101",
                     23115 => "11110000",
                     23116 => "01100110",
                     23117 => "10111101",
                     23118 => "11011000",
                     23119 => "00000011",
                     23120 => "11010000",
                     23121 => "01100001",
                     23122 => "00100000",
                     23123 => "01010100",
                     23124 => "11011100",
                     23125 => "11001010",
                     23126 => "00110000",
                     23127 => "01011011",
                     23128 => "10000110",
                     23129 => "00000001",
                     23130 => "10011000",
                     23131 => "01001000",
                     23132 => "10110101",
                     23133 => "00001111",
                     23134 => "11110000",
                     23135 => "01001100",
                     23136 => "10110101",
                     23137 => "00010110",
                     23138 => "11001001",
                     23139 => "00010101",
                     23140 => "10110000",
                     23141 => "01000110",
                     23142 => "11001001",
                     23143 => "00010001",
                     23144 => "11110000",
                     23145 => "01000010",
                     23146 => "11001001",
                     23147 => "00001101",
                     23148 => "11110000",
                     23149 => "00111110",
                     23150 => "10111101",
                     23151 => "11011000",
                     23152 => "00000011",
                     23153 => "11010000",
                     23154 => "00111001",
                     23155 => "10001010",
                     23156 => "00001010",
                     23157 => "00001010",
                     23158 => "00011000",
                     23159 => "01101001",
                     23160 => "00000100",
                     23161 => "10101010",
                     23162 => "00100000",
                     23163 => "00101111",
                     23164 => "11100011",
                     23165 => "10100110",
                     23166 => "00001000",
                     23167 => "10100100",
                     23168 => "00000001",
                     23169 => "10010000",
                     23170 => "00100000",
                     23171 => "10110101",
                     23172 => "00011110",
                     23173 => "00011001",
                     23174 => "00011110",
                     23175 => "00000000",
                     23176 => "00101001",
                     23177 => "10000000",
                     23178 => "11010000",
                     23179 => "00010001",
                     23180 => "10111001",
                     23181 => "10010001",
                     23182 => "00000100",
                     23183 => "00111101",
                     23184 => "00100111",
                     23185 => "11011010",
                     23186 => "11010000",
                     23187 => "00011000",
                     23188 => "10111001",
                     23189 => "10010001",
                     23190 => "00000100",
                     23191 => "00011101",
                     23192 => "00100111",
                     23193 => "11011010",
                     23194 => "10011001",
                     23195 => "10010001",
                     23196 => "00000100",
                     23197 => "00100000",
                     23198 => "10110110",
                     23199 => "11011010",
                     23200 => "01001100",
                     23201 => "10101100",
                     23202 => "11011010",
                     23203 => "10111001",
                     23204 => "10010001",
                     23205 => "00000100",
                     23206 => "00111101",
                     23207 => "00101110",
                     23208 => "11011010",
                     23209 => "10011001",
                     23210 => "10010001",
                     23211 => "00000100",
                     23212 => "01101000",
                     23213 => "10101000",
                     23214 => "10100110",
                     23215 => "00000001",
                     23216 => "11001010",
                     23217 => "00010000",
                     23218 => "10100101",
                     23219 => "10100110",
                     23220 => "00001000",
                     23221 => "01100000",
                     23222 => "10111001",
                     23223 => "00011110",
                     23224 => "00000000",
                     23225 => "00010101",
                     23226 => "00011110",
                     23227 => "00101001",
                     23228 => "00100000",
                     23229 => "11010000",
                     23230 => "00110011",
                     23231 => "10110101",
                     23232 => "00011110",
                     23233 => "11001001",
                     23234 => "00000110",
                     23235 => "10010000",
                     23236 => "00101110",
                     23237 => "10110101",
                     23238 => "00010110",
                     23239 => "11001001",
                     23240 => "00000101",
                     23241 => "11110000",
                     23242 => "00100111",
                     23243 => "10111001",
                     23244 => "00011110",
                     23245 => "00000000",
                     23246 => "00001010",
                     23247 => "10010000",
                     23248 => "00001010",
                     23249 => "10101001",
                     23250 => "00000110",
                     23251 => "00100000",
                     23252 => "00010011",
                     23253 => "11011010",
                     23254 => "00100000",
                     23255 => "10010101",
                     23256 => "11010111",
                     23257 => "10100100",
                     23258 => "00000001",
                     23259 => "10011000",
                     23260 => "10101010",
                     23261 => "00100000",
                     23262 => "10010101",
                     23263 => "11010111",
                     23264 => "10100110",
                     23265 => "00001000",
                     23266 => "10111101",
                     23267 => "00100101",
                     23268 => "00000001",
                     23269 => "00011000",
                     23270 => "01101001",
                     23271 => "00000100",
                     23272 => "10100110",
                     23273 => "00000001",
                     23274 => "00100000",
                     23275 => "00010011",
                     23276 => "11011010",
                     23277 => "10100110",
                     23278 => "00001000",
                     23279 => "11111110",
                     23280 => "00100101",
                     23281 => "00000001",
                     23282 => "01100000",
                     23283 => "10111001",
                     23284 => "00011110",
                     23285 => "00000000",
                     23286 => "11001001",
                     23287 => "00000110",
                     23288 => "10010000",
                     23289 => "00011101",
                     23290 => "10111001",
                     23291 => "00010110",
                     23292 => "00000000",
                     23293 => "11001001",
                     23294 => "00000101",
                     23295 => "11110000",
                     23296 => "11110001",
                     23297 => "00100000",
                     23298 => "10010101",
                     23299 => "11010111",
                     23300 => "10100100",
                     23301 => "00000001",
                     23302 => "10111001",
                     23303 => "00100101",
                     23304 => "00000001",
                     23305 => "00011000",
                     23306 => "01101001",
                     23307 => "00000100",
                     23308 => "10100110",
                     23309 => "00001000",
                     23310 => "00100000",
                     23311 => "00010011",
                     23312 => "11011010",
                     23313 => "10100110",
                     23314 => "00000001",
                     23315 => "11111110",
                     23316 => "00100101",
                     23317 => "00000001",
                     23318 => "01100000",
                     23319 => "10011000",
                     23320 => "10101010",
                     23321 => "00100000",
                     23322 => "00011110",
                     23323 => "11011011",
                     23324 => "10100110",
                     23325 => "00001000",
                     23326 => "10110101",
                     23327 => "00010110",
                     23328 => "11001001",
                     23329 => "00001101",
                     23330 => "11110000",
                     23331 => "00100010",
                     23332 => "11001001",
                     23333 => "00010001",
                     23334 => "11110000",
                     23335 => "00011110",
                     23336 => "11001001",
                     23337 => "00000101",
                     23338 => "11110000",
                     23339 => "00011010",
                     23340 => "11001001",
                     23341 => "00010010",
                     23342 => "11110000",
                     23343 => "00001000",
                     23344 => "11001001",
                     23345 => "00001110",
                     23346 => "11110000",
                     23347 => "00000100",
                     23348 => "11001001",
                     23349 => "00000111",
                     23350 => "10110000",
                     23351 => "00001110",
                     23352 => "10110101",
                     23353 => "01011000",
                     23354 => "01001001",
                     23355 => "11111111",
                     23356 => "10101000",
                     23357 => "11001000",
                     23358 => "10010100",
                     23359 => "01011000",
                     23360 => "10110101",
                     23361 => "01000110",
                     23362 => "01001001",
                     23363 => "00000011",
                     23364 => "10010101",
                     23365 => "01000110",
                     23366 => "01100000",
                     23367 => "10101001",
                     23368 => "11111111",
                     23369 => "10011101",
                     23370 => "10100010",
                     23371 => "00000011",
                     23372 => "10101101",
                     23373 => "01000111",
                     23374 => "00000111",
                     23375 => "11010000",
                     23376 => "00101001",
                     23377 => "10110101",
                     23378 => "00011110",
                     23379 => "00110000",
                     23380 => "00100101",
                     23381 => "10110101",
                     23382 => "00010110",
                     23383 => "11001001",
                     23384 => "00100100",
                     23385 => "11010000",
                     23386 => "00000110",
                     23387 => "10110101",
                     23388 => "00011110",
                     23389 => "10101010",
                     23390 => "00100000",
                     23391 => "01100001",
                     23392 => "11011011",
                     23393 => "00100000",
                     23394 => "01000011",
                     23395 => "11011100",
                     23396 => "10110000",
                     23397 => "00010100",
                     23398 => "10001010",
                     23399 => "00100000",
                     23400 => "01010110",
                     23401 => "11011100",
                     23402 => "10110101",
                     23403 => "11001111",
                     23404 => "10000101",
                     23405 => "00000000",
                     23406 => "10001010",
                     23407 => "01001000",
                     23408 => "00100000",
                     23409 => "00101101",
                     23410 => "11100011",
                     23411 => "01101000",
                     23412 => "10101010",
                     23413 => "10010000",
                     23414 => "00000011",
                     23415 => "00100000",
                     23416 => "10111110",
                     23417 => "11011011",
                     23418 => "10100110",
                     23419 => "00001000",
                     23420 => "01100000",
                     23421 => "10101101",
                     23422 => "01000111",
                     23423 => "00000111",
                     23424 => "11010000",
                     23425 => "00110111",
                     23426 => "10011101",
                     23427 => "10100010",
                     23428 => "00000011",
                     23429 => "00100000",
                     23430 => "01000011",
                     23431 => "11011100",
                     23432 => "10110000",
                     23433 => "00101111",
                     23434 => "10101001",
                     23435 => "00000010",
                     23436 => "10000101",
                     23437 => "00000000",
                     23438 => "10100110",
                     23439 => "00001000",
                     23440 => "00100000",
                     23441 => "01010100",
                     23442 => "11011100",
                     23443 => "00101001",
                     23444 => "00000010",
                     23445 => "11010000",
                     23446 => "00100010",
                     23447 => "10111001",
                     23448 => "10101101",
                     23449 => "00000100",
                     23450 => "11001001",
                     23451 => "00100000",
                     23452 => "10010000",
                     23453 => "00000101",
                     23454 => "00100000",
                     23455 => "00101101",
                     23456 => "11100011",
                     23457 => "10110000",
                     23458 => "00011001",
                     23459 => "10111001",
                     23460 => "10101101",
                     23461 => "00000100",
                     23462 => "00011000",
                     23463 => "01101001",
                     23464 => "10000000",
                     23465 => "10011001",
                     23466 => "10101101",
                     23467 => "00000100",
                     23468 => "10111001",
                     23469 => "10101111",
                     23470 => "00000100",
                     23471 => "00011000",
                     23472 => "01101001",
                     23473 => "10000000",
                     23474 => "10011001",
                     23475 => "10101111",
                     23476 => "00000100",
                     23477 => "11000110",
                     23478 => "00000000",
                     23479 => "11010000",
                     23480 => "11010101",
                     23481 => "10100110",
                     23482 => "00001000",
                     23483 => "01100000",
                     23484 => "10100110",
                     23485 => "00001000",
                     23486 => "10111001",
                     23487 => "10101111",
                     23488 => "00000100",
                     23489 => "00111000",
                     23490 => "11101101",
                     23491 => "10101101",
                     23492 => "00000100",
                     23493 => "11001001",
                     23494 => "00000100",
                     23495 => "10110000",
                     23496 => "00001000",
                     23497 => "10100101",
                     23498 => "10011111",
                     23499 => "00010000",
                     23500 => "00000100",
                     23501 => "10101001",
                     23502 => "00000001",
                     23503 => "10000101",
                     23504 => "10011111",
                     23505 => "10101101",
                     23506 => "10101111",
                     23507 => "00000100",
                     23508 => "00111000",
                     23509 => "11111001",
                     23510 => "10101101",
                     23511 => "00000100",
                     23512 => "11001001",
                     23513 => "00000110",
                     23514 => "10110000",
                     23515 => "00011011",
                     23516 => "10100101",
                     23517 => "10011111",
                     23518 => "00110000",
                     23519 => "00010111",
                     23520 => "10100101",
                     23521 => "00000000",
                     23522 => "10110100",
                     23523 => "00010110",
                     23524 => "11000000",
                     23525 => "00101011",
                     23526 => "11110000",
                     23527 => "00000101",
                     23528 => "11000000",
                     23529 => "00101100",
                     23530 => "11110000",
                     23531 => "00000001",
                     23532 => "10001010",
                     23533 => "10100110",
                     23534 => "00001000",
                     23535 => "10011101",
                     23536 => "10100010",
                     23537 => "00000011",
                     23538 => "10101001",
                     23539 => "00000000",
                     23540 => "10000101",
                     23541 => "00011101",
                     23542 => "01100000",
                     23543 => "10101001",
                     23544 => "00000001",
                     23545 => "10000101",
                     23546 => "00000000",
                     23547 => "10101101",
                     23548 => "10101110",
                     23549 => "00000100",
                     23550 => "00111000",
                     23551 => "11111001",
                     23552 => "10101100",
                     23553 => "00000100",
                     23554 => "11001001",
                     23555 => "00001000",
                     23556 => "10010000",
                     23557 => "00001101",
                     23558 => "11100110",
                     23559 => "00000000",
                     23560 => "10111001",
                     23561 => "10101110",
                     23562 => "00000100",
                     23563 => "00011000",
                     23564 => "11101101",
                     23565 => "10101100",
                     23566 => "00000100",
                     23567 => "11001001",
                     23568 => "00001001",
                     23569 => "10110000",
                     23570 => "00000011",
                     23571 => "00100000",
                     23572 => "01010011",
                     23573 => "11011111",
                     23574 => "10100110",
                     23575 => "00001000",
                     23576 => "01100000",
                     23577 => "10000000",
                     23578 => "00000000",
                     23579 => "10101000",
                     23580 => "10110101",
                     23581 => "11001111",
                     23582 => "00011000",
                     23583 => "01111001",
                     23584 => "00011000",
                     23585 => "11011100",
                     23586 => "00101100",
                     23587 => "10110101",
                     23588 => "11001111",
                     23589 => "10100100",
                     23590 => "00001110",
                     23591 => "11000000",
                     23592 => "00001011",
                     23593 => "11110000",
                     23594 => "00010111",
                     23595 => "10110100",
                     23596 => "10110110",
                     23597 => "11000000",
                     23598 => "00000001",
                     23599 => "11010000",
                     23600 => "00010001",
                     23601 => "00111000",
                     23602 => "11101001",
                     23603 => "00100000",
                     23604 => "10000101",
                     23605 => "11001110",
                     23606 => "10011000",
                     23607 => "11101001",
                     23608 => "00000000",
                     23609 => "10000101",
                     23610 => "10110101",
                     23611 => "10101001",
                     23612 => "00000000",
                     23613 => "10000101",
                     23614 => "10011111",
                     23615 => "10001101",
                     23616 => "00110011",
                     23617 => "00000100",
                     23618 => "01100000",
                     23619 => "10101101",
                     23620 => "11010000",
                     23621 => "00000011",
                     23622 => "11001001",
                     23623 => "11110000",
                     23624 => "10110000",
                     23625 => "00001001",
                     23626 => "10100100",
                     23627 => "10110101",
                     23628 => "10001000",
                     23629 => "11010000",
                     23630 => "00000100",
                     23631 => "10100101",
                     23632 => "11001110",
                     23633 => "11001001",
                     23634 => "11010000",
                     23635 => "01100000",
                     23636 => "10100101",
                     23637 => "00001000",
                     23638 => "00001010",
                     23639 => "00001010",
                     23640 => "00011000",
                     23641 => "01101001",
                     23642 => "00000100",
                     23643 => "10101000",
                     23644 => "10101101",
                     23645 => "11010001",
                     23646 => "00000011",
                     23647 => "00101001",
                     23648 => "00001111",
                     23649 => "11001001",
                     23650 => "00001111",
                     23651 => "01100000",
                     23652 => "00100000",
                     23653 => "00010000",
                     23654 => "10101101",
                     23655 => "00010110",
                     23656 => "00000111",
                     23657 => "11010000",
                     23658 => "00101110",
                     23659 => "10100101",
                     23660 => "00001110",
                     23661 => "11001001",
                     23662 => "00001011",
                     23663 => "11110000",
                     23664 => "00101000",
                     23665 => "11001001",
                     23666 => "00000100",
                     23667 => "10010000",
                     23668 => "00100100",
                     23669 => "10101001",
                     23670 => "00000001",
                     23671 => "10101100",
                     23672 => "00000100",
                     23673 => "00000111",
                     23674 => "11010000",
                     23675 => "00001010",
                     23676 => "10100101",
                     23677 => "00011101",
                     23678 => "11110000",
                     23679 => "00000100",
                     23680 => "11001001",
                     23681 => "00000011",
                     23682 => "11010000",
                     23683 => "00000100",
                     23684 => "10101001",
                     23685 => "00000010",
                     23686 => "10000101",
                     23687 => "00011101",
                     23688 => "10100101",
                     23689 => "10110101",
                     23690 => "11001001",
                     23691 => "00000001",
                     23692 => "11010000",
                     23693 => "00001011",
                     23694 => "10101001",
                     23695 => "11111111",
                     23696 => "10001101",
                     23697 => "10010000",
                     23698 => "00000100",
                     23699 => "10100101",
                     23700 => "11001110",
                     23701 => "11001001",
                     23702 => "11001111",
                     23703 => "10010000",
                     23704 => "00000001",
                     23705 => "01100000",
                     23706 => "10100000",
                     23707 => "00000010",
                     23708 => "10101101",
                     23709 => "00010100",
                     23710 => "00000111",
                     23711 => "11010000",
                     23712 => "00001100",
                     23713 => "10101101",
                     23714 => "01010100",
                     23715 => "00000111",
                     23716 => "11010000",
                     23717 => "00000111",
                     23718 => "10001000",
                     23719 => "10101101",
                     23720 => "00000100",
                     23721 => "00000111",
                     23722 => "11010000",
                     23723 => "00000001",
                     23724 => "10001000",
                     23725 => "10111001",
                     23726 => "10110101",
                     23727 => "11100011",
                     23728 => "10000101",
                     23729 => "11101011",
                     23730 => "10101000",
                     23731 => "10101110",
                     23732 => "01010100",
                     23733 => "00000111",
                     23734 => "10101101",
                     23735 => "00010100",
                     23736 => "00000111",
                     23737 => "11110000",
                     23738 => "00000001",
                     23739 => "11101000",
                     23740 => "10100101",
                     23741 => "11001110",
                     23742 => "11011101",
                     23743 => "01100100",
                     23744 => "11011100",
                     23745 => "10010000",
                     23746 => "00111011",
                     23747 => "00100000",
                     23748 => "11110001",
                     23749 => "11100011",
                     23750 => "11110000",
                     23751 => "00110110",
                     23752 => "00100000",
                     23753 => "10101001",
                     23754 => "11011111",
                     23755 => "10110000",
                     23756 => "01010101",
                     23757 => "10100100",
                     23758 => "10011111",
                     23759 => "00010000",
                     23760 => "00101101",
                     23761 => "10100100",
                     23762 => "00000100",
                     23763 => "11000000",
                     23764 => "00000100",
                     23765 => "10010000",
                     23766 => "00100111",
                     23767 => "00100000",
                     23768 => "10010111",
                     23769 => "11011111",
                     23770 => "10110000",
                     23771 => "00010000",
                     23772 => "10101100",
                     23773 => "01001110",
                     23774 => "00000111",
                     23775 => "11110000",
                     23776 => "00010011",
                     23777 => "10101100",
                     23778 => "10000100",
                     23779 => "00000111",
                     23780 => "11010000",
                     23781 => "00001110",
                     23782 => "00100000",
                     23783 => "11110010",
                     23784 => "10111100",
                     23785 => "01001100",
                     23786 => "11111110",
                     23787 => "11011100",
                     23788 => "11001001",
                     23789 => "00100110",
                     23790 => "11110000",
                     23791 => "00000100",
                     23792 => "10101001",
                     23793 => "00000010",
                     23794 => "10000101",
                     23795 => "11111111",
                     23796 => "10100000",
                     23797 => "00000001",
                     23798 => "10101101",
                     23799 => "01001110",
                     23800 => "00000111",
                     23801 => "11010000",
                     23802 => "00000001",
                     23803 => "10001000",
                     23804 => "10000100",
                     23805 => "10011111",
                     23806 => "10100100",
                     23807 => "11101011",
                     23808 => "10100101",
                     23809 => "11001110",
                     23810 => "11001001",
                     23811 => "11001111",
                     23812 => "10110000",
                     23813 => "01100000",
                     23814 => "00100000",
                     23815 => "11110000",
                     23816 => "11100011",
                     23817 => "00100000",
                     23818 => "10101001",
                     23819 => "11011111",
                     23820 => "10110000",
                     23821 => "00010100",
                     23822 => "01001000",
                     23823 => "00100000",
                     23824 => "11110000",
                     23825 => "11100011",
                     23826 => "10000101",
                     23827 => "00000000",
                     23828 => "01101000",
                     23829 => "10000101",
                     23830 => "00000001",
                     23831 => "11010000",
                     23832 => "00001100",
                     23833 => "10100101",
                     23834 => "00000000",
                     23835 => "11110000",
                     23836 => "01001001",
                     23837 => "00100000",
                     23838 => "10101001",
                     23839 => "11011111",
                     23840 => "10010000",
                     23841 => "00000011",
                     23842 => "01001100",
                     23843 => "00001101",
                     23844 => "11011110",
                     23845 => "00100000",
                     23846 => "10100010",
                     23847 => "11011111",
                     23848 => "10110000",
                     23849 => "00111100",
                     23850 => "10100100",
                     23851 => "10011111",
                     23852 => "00110000",
                     23853 => "00111000",
                     23854 => "11001001",
                     23855 => "11000101",
                     23856 => "11010000",
                     23857 => "00000011",
                     23858 => "01001100",
                     23859 => "00010110",
                     23860 => "11011110",
                     23861 => "00100000",
                     23862 => "11000101",
                     23863 => "11011110",
                     23864 => "11110000",
                     23865 => "00101100",
                     23866 => "10101100",
                     23867 => "00001110",
                     23868 => "00000111",
                     23869 => "11010000",
                     23870 => "00100011",
                     23871 => "10100100",
                     23872 => "00000100",
                     23873 => "11000000",
                     23874 => "00000110",
                     23875 => "10010000",
                     23876 => "00000111",
                     23877 => "10100101",
                     23878 => "01000101",
                     23879 => "10000101",
                     23880 => "00000000",
                     23881 => "01001100",
                     23882 => "01010011",
                     23883 => "11011111",
                     23884 => "00100000",
                     23885 => "11001100",
                     23886 => "11011110",
                     23887 => "10101001",
                     23888 => "11110000",
                     23889 => "00100101",
                     23890 => "11001110",
                     23891 => "10000101",
                     23892 => "11001110",
                     23893 => "00100000",
                     23894 => "11110000",
                     23895 => "11011110",
                     23896 => "10101001",
                     23897 => "00000000",
                     23898 => "10000101",
                     23899 => "10011111",
                     23900 => "10001101",
                     23901 => "00110011",
                     23902 => "00000100",
                     23903 => "10001101",
                     23904 => "10000100",
                     23905 => "00000100",
                     23906 => "10101001",
                     23907 => "00000000",
                     23908 => "10000101",
                     23909 => "00011101",
                     23910 => "10100100",
                     23911 => "11101011",
                     23912 => "11001000",
                     23913 => "11001000",
                     23914 => "10101001",
                     23915 => "00000010",
                     23916 => "10000101",
                     23917 => "00000000",
                     23918 => "11001000",
                     23919 => "10000100",
                     23920 => "11101011",
                     23921 => "10100101",
                     23922 => "11001110",
                     23923 => "11001001",
                     23924 => "00100000",
                     23925 => "10010000",
                     23926 => "00010110",
                     23927 => "11001001",
                     23928 => "11100100",
                     23929 => "10110000",
                     23930 => "00101000",
                     23931 => "00100000",
                     23932 => "11110100",
                     23933 => "11100011",
                     23934 => "11110000",
                     23935 => "00001101",
                     23936 => "11001001",
                     23937 => "00011100",
                     23938 => "11110000",
                     23939 => "00001001",
                     23940 => "11001001",
                     23941 => "01101011",
                     23942 => "11110000",
                     23943 => "00000101",
                     23944 => "00100000",
                     23945 => "10100010",
                     23946 => "11011111",
                     23947 => "10010000",
                     23948 => "00010111",
                     23949 => "10100100",
                     23950 => "11101011",
                     23951 => "11001000",
                     23952 => "10100101",
                     23953 => "11001110",
                     23954 => "11001001",
                     23955 => "00001000",
                     23956 => "10010000",
                     23957 => "00001101",
                     23958 => "11001001",
                     23959 => "11010000",
                     23960 => "10110000",
                     23961 => "00001001",
                     23962 => "00100000",
                     23963 => "11110100",
                     23964 => "11100011",
                     23965 => "11010000",
                     23966 => "00000101",
                     23967 => "11000110",
                     23968 => "00000000",
                     23969 => "11010000",
                     23970 => "11001011",
                     23971 => "01100000",
                     23972 => "00100000",
                     23973 => "11000101",
                     23974 => "11011110",
                     23975 => "11110000",
                     23976 => "01100001",
                     23977 => "00100000",
                     23978 => "10100010",
                     23979 => "11011111",
                     23980 => "10010000",
                     23981 => "00000011",
                     23982 => "01001100",
                     23983 => "00110110",
                     23984 => "11011110",
                     23985 => "00100000",
                     23986 => "10101001",
                     23987 => "11011111",
                     23988 => "10110000",
                     23989 => "01010111",
                     23990 => "00100000",
                     23991 => "11100101",
                     23992 => "11011110",
                     23993 => "10010000",
                     23994 => "00001000",
                     23995 => "10101101",
                     23996 => "00001110",
                     23997 => "00000111",
                     23998 => "11010000",
                     23999 => "01001010",
                     24000 => "01001100",
                     24001 => "00000111",
                     24002 => "11011110",
                     24003 => "10100100",
                     24004 => "00011101",
                     24005 => "11000000",
                     24006 => "00000000",
                     24007 => "11010000",
                     24008 => "00111110",
                     24009 => "10100100",
                     24010 => "00110011",
                     24011 => "10001000",
                     24012 => "11010000",
                     24013 => "00111001",
                     24014 => "11001001",
                     24015 => "01101100",
                     24016 => "11110000",
                     24017 => "00000100",
                     24018 => "11001001",
                     24019 => "00011111",
                     24020 => "11010000",
                     24021 => "00110001",
                     24022 => "10101101",
                     24023 => "11000100",
                     24024 => "00000011",
                     24025 => "11010000",
                     24026 => "00000100",
                     24027 => "10100000",
                     24028 => "00010000",
                     24029 => "10000100",
                     24030 => "11111111",
                     24031 => "00001001",
                     24032 => "00100000",
                     24033 => "10001101",
                     24034 => "11000100",
                     24035 => "00000011",
                     24036 => "10100101",
                     24037 => "10000110",
                     24038 => "00101001",
                     24039 => "00001111",
                     24040 => "11110000",
                     24041 => "00001110",
                     24042 => "10100000",
                     24043 => "00000000",
                     24044 => "10101101",
                     24045 => "00011010",
                     24046 => "00000111",
                     24047 => "11110000",
                     24048 => "00000001",
                     24049 => "11001000",
                     24050 => "10111001",
                     24051 => "00001011",
                     24052 => "11011110",
                     24053 => "10001101",
                     24054 => "11011110",
                     24055 => "00000110",
                     24056 => "10100101",
                     24057 => "00001110",
                     24058 => "11001001",
                     24059 => "00000111",
                     24060 => "11110000",
                     24061 => "00001100",
                     24062 => "11001001",
                     24063 => "00001000",
                     24064 => "11010000",
                     24065 => "00001000",
                     24066 => "10101001",
                     24067 => "00000010",
                     24068 => "10000101",
                     24069 => "00001110",
                     24070 => "01100000",
                     24071 => "00100000",
                     24072 => "01010011",
                     24073 => "11011111",
                     24074 => "01100000",
                     24075 => "10000101",
                     24076 => "00101011",
                     24077 => "00100000",
                     24078 => "00100100",
                     24079 => "11011110",
                     24080 => "11101110",
                     24081 => "01001000",
                     24082 => "00000111",
                     24083 => "01001100",
                     24084 => "00000011",
                     24085 => "10111100",
                     24086 => "10101001",
                     24087 => "00000000",
                     24088 => "10001101",
                     24089 => "01110010",
                     24090 => "00000111",
                     24091 => "10101001",
                     24092 => "00000010",
                     24093 => "10001101",
                     24094 => "01110000",
                     24095 => "00000111",
                     24096 => "10101001",
                     24097 => "00011000",
                     24098 => "10000101",
                     24099 => "01010111",
                     24100 => "10100100",
                     24101 => "00000010",
                     24102 => "10101001",
                     24103 => "00000000",
                     24104 => "10010001",
                     24105 => "00000110",
                     24106 => "01001100",
                     24107 => "01001101",
                     24108 => "10001010",
                     24109 => "11111001",
                     24110 => "00000111",
                     24111 => "11111111",
                     24112 => "00000000",
                     24113 => "00011000",
                     24114 => "00100010",
                     24115 => "01010000",
                     24116 => "01101000",
                     24117 => "10010000",
                     24118 => "10100100",
                     24119 => "00000100",
                     24120 => "11000000",
                     24121 => "00000110",
                     24122 => "10010000",
                     24123 => "00000100",
                     24124 => "11000000",
                     24125 => "00001010",
                     24126 => "10010000",
                     24127 => "00000001",
                     24128 => "01100000",
                     24129 => "11001001",
                     24130 => "00100100",
                     24131 => "11110000",
                     24132 => "00000100",
                     24133 => "11001001",
                     24134 => "00100101",
                     24135 => "11010000",
                     24136 => "00111001",
                     24137 => "10100101",
                     24138 => "00001110",
                     24139 => "11001001",
                     24140 => "00000101",
                     24141 => "11110000",
                     24142 => "01000001",
                     24143 => "10101001",
                     24144 => "00000001",
                     24145 => "10000101",
                     24146 => "00110011",
                     24147 => "11101110",
                     24148 => "00100011",
                     24149 => "00000111",
                     24150 => "10100101",
                     24151 => "00001110",
                     24152 => "11001001",
                     24153 => "00000100",
                     24154 => "11110000",
                     24155 => "00011111",
                     24156 => "10101001",
                     24157 => "00110011",
                     24158 => "00100000",
                     24159 => "00010110",
                     24160 => "10010111",
                     24161 => "10101001",
                     24162 => "10000000",
                     24163 => "10000101",
                     24164 => "11111100",
                     24165 => "01001010",
                     24166 => "10001101",
                     24167 => "00010011",
                     24168 => "00000111",
                     24169 => "10100010",
                     24170 => "00000100",
                     24171 => "10100101",
                     24172 => "11001110",
                     24173 => "10001101",
                     24174 => "00001111",
                     24175 => "00000111",
                     24176 => "11011101",
                     24177 => "00110001",
                     24178 => "11011110",
                     24179 => "10110000",
                     24180 => "00000011",
                     24181 => "11001010",
                     24182 => "11010000",
                     24183 => "11111000",
                     24184 => "10001110",
                     24185 => "00001111",
                     24186 => "00000001",
                     24187 => "10101001",
                     24188 => "00000100",
                     24189 => "10000101",
                     24190 => "00001110",
                     24191 => "01001100",
                     24192 => "10010000",
                     24193 => "11011110",
                     24194 => "11001001",
                     24195 => "00100110",
                     24196 => "11010000",
                     24197 => "00001010",
                     24198 => "10100101",
                     24199 => "11001110",
                     24200 => "11001001",
                     24201 => "00100000",
                     24202 => "10110000",
                     24203 => "00000100",
                     24204 => "10101001",
                     24205 => "00000001",
                     24206 => "10000101",
                     24207 => "00001110",
                     24208 => "10101001",
                     24209 => "00000011",
                     24210 => "10000101",
                     24211 => "00011101",
                     24212 => "10101001",
                     24213 => "00000000",
                     24214 => "10000101",
                     24215 => "01010111",
                     24216 => "10001101",
                     24217 => "00000101",
                     24218 => "00000111",
                     24219 => "10100101",
                     24220 => "10000110",
                     24221 => "00111000",
                     24222 => "11101101",
                     24223 => "00011100",
                     24224 => "00000111",
                     24225 => "11001001",
                     24226 => "00010000",
                     24227 => "10110000",
                     24228 => "00000100",
                     24229 => "10101001",
                     24230 => "00000010",
                     24231 => "10000101",
                     24232 => "00110011",
                     24233 => "10100100",
                     24234 => "00110011",
                     24235 => "10100101",
                     24236 => "00000110",
                     24237 => "00001010",
                     24238 => "00001010",
                     24239 => "00001010",
                     24240 => "00001010",
                     24241 => "00011000",
                     24242 => "01111001",
                     24243 => "00101100",
                     24244 => "11011110",
                     24245 => "10000101",
                     24246 => "10000110",
                     24247 => "10100101",
                     24248 => "00000110",
                     24249 => "11010000",
                     24250 => "00001001",
                     24251 => "10101101",
                     24252 => "00011011",
                     24253 => "00000111",
                     24254 => "00011000",
                     24255 => "01111001",
                     24256 => "00101110",
                     24257 => "11011110",
                     24258 => "10000101",
                     24259 => "01101101",
                     24260 => "01100000",
                     24261 => "11001001",
                     24262 => "01011111",
                     24263 => "11110000",
                     24264 => "00000010",
                     24265 => "11001001",
                     24266 => "01100000",
                     24267 => "01100000",
                     24268 => "00100000",
                     24269 => "11100101",
                     24270 => "11011110",
                     24271 => "10010000",
                     24272 => "00010011",
                     24273 => "10101001",
                     24274 => "01110000",
                     24275 => "10001101",
                     24276 => "00001001",
                     24277 => "00000111",
                     24278 => "10101001",
                     24279 => "11111000",
                     24280 => "10001101",
                     24281 => "11011011",
                     24282 => "00000110",
                     24283 => "10101001",
                     24284 => "00000011",
                     24285 => "10001101",
                     24286 => "10000110",
                     24287 => "00000111",
                     24288 => "01001010",
                     24289 => "10001101",
                     24290 => "00001110",
                     24291 => "00000111",
                     24292 => "01100000",
                     24293 => "11001001",
                     24294 => "01100111",
                     24295 => "11110000",
                     24296 => "00000101",
                     24297 => "11001001",
                     24298 => "01101000",
                     24299 => "00011000",
                     24300 => "11010000",
                     24301 => "00000001",
                     24302 => "00111000",
                     24303 => "01100000",
                     24304 => "10100101",
                     24305 => "00001011",
                     24306 => "00101001",
                     24307 => "00000100",
                     24308 => "11110000",
                     24309 => "01011100",
                     24310 => "10100101",
                     24311 => "00000000",
                     24312 => "11001001",
                     24313 => "00010001",
                     24314 => "11010000",
                     24315 => "01010110",
                     24316 => "10100101",
                     24317 => "00000001",
                     24318 => "11001001",
                     24319 => "00010000",
                     24320 => "11010000",
                     24321 => "01010000",
                     24322 => "10101001",
                     24323 => "00101000",
                     24324 => "10001101",
                     24325 => "11011110",
                     24326 => "00000110",
                     24327 => "10101001",
                     24328 => "00000011",
                     24329 => "10000101",
                     24330 => "00001110",
                     24331 => "10101001",
                     24332 => "00010000",
                     24333 => "10000101",
                     24334 => "11111111",
                     24335 => "10101001",
                     24336 => "00100000",
                     24337 => "10001101",
                     24338 => "11000100",
                     24339 => "00000011",
                     24340 => "10101101",
                     24341 => "11010110",
                     24342 => "00000110",
                     24343 => "11110000",
                     24344 => "00111001",
                     24345 => "00101001",
                     24346 => "00000011",
                     24347 => "00001010",
                     24348 => "00001010",
                     24349 => "10101010",
                     24350 => "10100101",
                     24351 => "10000110",
                     24352 => "11001001",
                     24353 => "01100000",
                     24354 => "10010000",
                     24355 => "00000110",
                     24356 => "11101000",
                     24357 => "11001001",
                     24358 => "10100000",
                     24359 => "10010000",
                     24360 => "00000001",
                     24361 => "11101000",
                     24362 => "10111100",
                     24363 => "11110010",
                     24364 => "10000111",
                     24365 => "10001000",
                     24366 => "10001100",
                     24367 => "01011111",
                     24368 => "00000111",
                     24369 => "10111110",
                     24370 => "10110100",
                     24371 => "10011100",
                     24372 => "10111101",
                     24373 => "10111100",
                     24374 => "10011100",
                     24375 => "10001101",
                     24376 => "01010000",
                     24377 => "00000111",
                     24378 => "10101001",
                     24379 => "10000000",
                     24380 => "10000101",
                     24381 => "11111100",
                     24382 => "10101001",
                     24383 => "00000000",
                     24384 => "10001101",
                     24385 => "01010001",
                     24386 => "00000111",
                     24387 => "10001101",
                     24388 => "01100000",
                     24389 => "00000111",
                     24390 => "10001101",
                     24391 => "01011100",
                     24392 => "00000111",
                     24393 => "10001101",
                     24394 => "01010010",
                     24395 => "00000111",
                     24396 => "11101110",
                     24397 => "01011101",
                     24398 => "00000111",
                     24399 => "11101110",
                     24400 => "01010111",
                     24401 => "00000111",
                     24402 => "01100000",
                     24403 => "10101001",
                     24404 => "00000000",
                     24405 => "10100100",
                     24406 => "01010111",
                     24407 => "10100110",
                     24408 => "00000000",
                     24409 => "11001010",
                     24410 => "11010000",
                     24411 => "00001010",
                     24412 => "11101000",
                     24413 => "11000000",
                     24414 => "00000000",
                     24415 => "00110000",
                     24416 => "00101000",
                     24417 => "10101001",
                     24418 => "11111111",
                     24419 => "01001100",
                     24420 => "01101110",
                     24421 => "11011111",
                     24422 => "10100010",
                     24423 => "00000010",
                     24424 => "11000000",
                     24425 => "00000001",
                     24426 => "00010000",
                     24427 => "00011101",
                     24428 => "10101001",
                     24429 => "00000001",
                     24430 => "10100000",
                     24431 => "00010000",
                     24432 => "10001100",
                     24433 => "10000101",
                     24434 => "00000111",
                     24435 => "10100000",
                     24436 => "00000000",
                     24437 => "10000100",
                     24438 => "01010111",
                     24439 => "11001001",
                     24440 => "00000000",
                     24441 => "00010000",
                     24442 => "00000001",
                     24443 => "10001000",
                     24444 => "10000100",
                     24445 => "00000000",
                     24446 => "00011000",
                     24447 => "01100101",
                     24448 => "10000110",
                     24449 => "10000101",
                     24450 => "10000110",
                     24451 => "10100101",
                     24452 => "01101101",
                     24453 => "01100101",
                     24454 => "00000000",
                     24455 => "10000101",
                     24456 => "01101101",
                     24457 => "10001010",
                     24458 => "01001001",
                     24459 => "11111111",
                     24460 => "00101101",
                     24461 => "10010000",
                     24462 => "00000100",
                     24463 => "10001101",
                     24464 => "10010000",
                     24465 => "00000100",
                     24466 => "01100000",
                     24467 => "00010000",
                     24468 => "01100001",
                     24469 => "10001000",
                     24470 => "11000100",
                     24471 => "00100000",
                     24472 => "10111000",
                     24473 => "11011111",
                     24474 => "11011101",
                     24475 => "10010011",
                     24476 => "11011111",
                     24477 => "01100000",
                     24478 => "00100100",
                     24479 => "01101101",
                     24480 => "10001010",
                     24481 => "11000110",
                     24482 => "00100000",
                     24483 => "10111000",
                     24484 => "11011111",
                     24485 => "11011101",
                     24486 => "10011110",
                     24487 => "11011111",
                     24488 => "01100000",
                     24489 => "11001001",
                     24490 => "11000010",
                     24491 => "11110000",
                     24492 => "00000110",
                     24493 => "11001001",
                     24494 => "11000011",
                     24495 => "11110000",
                     24496 => "00000010",
                     24497 => "00011000",
                     24498 => "01100000",
                     24499 => "10101001",
                     24500 => "00000001",
                     24501 => "10000101",
                     24502 => "11111110",
                     24503 => "01100000",
                     24504 => "10101000",
                     24505 => "00101001",
                     24506 => "11000000",
                     24507 => "00001010",
                     24508 => "00101010",
                     24509 => "00101010",
                     24510 => "10101010",
                     24511 => "10011000",
                     24512 => "01100000",
                     24513 => "00000001",
                     24514 => "00000001",
                     24515 => "00000010",
                     24516 => "00000010",
                     24517 => "00000010",
                     24518 => "00000101",
                     24519 => "00010000",
                     24520 => "11110000",
                     24521 => "10110101",
                     24522 => "00011110",
                     24523 => "00101001",
                     24524 => "00100000",
                     24525 => "11010000",
                     24526 => "11110001",
                     24527 => "00100000",
                     24528 => "01100011",
                     24529 => "11100001",
                     24530 => "10010000",
                     24531 => "11101100",
                     24532 => "10110100",
                     24533 => "00010110",
                     24534 => "11000000",
                     24535 => "00010010",
                     24536 => "11010000",
                     24537 => "00000110",
                     24538 => "10110101",
                     24539 => "11001111",
                     24540 => "11001001",
                     24541 => "00100101",
                     24542 => "10010000",
                     24543 => "11100000",
                     24544 => "11000000",
                     24545 => "00001110",
                     24546 => "11010000",
                     24547 => "00000011",
                     24548 => "01001100",
                     24549 => "01101011",
                     24550 => "11100001",
                     24551 => "11000000",
                     24552 => "00000101",
                     24553 => "11010000",
                     24554 => "00000011",
                     24555 => "01001100",
                     24556 => "10001101",
                     24557 => "11100001",
                     24558 => "11000000",
                     24559 => "00010010",
                     24560 => "11110000",
                     24561 => "00001000",
                     24562 => "11000000",
                     24563 => "00101110",
                     24564 => "11110000",
                     24565 => "00000100",
                     24566 => "11000000",
                     24567 => "00000111",
                     24568 => "10110000",
                     24569 => "01110100",
                     24570 => "00100000",
                     24571 => "10110110",
                     24572 => "11100001",
                     24573 => "11010000",
                     24574 => "00000011",
                     24575 => "01001100",
                     24576 => "11101010",
                     24577 => "11100000",
                     24578 => "00100000",
                     24579 => "10111101",
                     24580 => "11100001",
                     24581 => "11110000",
                     24582 => "11111000",
                     24583 => "11001001",
                     24584 => "00100011",
                     24585 => "11010000",
                     24586 => "01100100",
                     24587 => "10100100",
                     24588 => "00000010",
                     24589 => "10101001",
                     24590 => "00000000",
                     24591 => "10010001",
                     24592 => "00000110",
                     24593 => "10110101",
                     24594 => "00010110",
                     24595 => "11001001",
                     24596 => "00010101",
                     24597 => "10110000",
                     24598 => "00001100",
                     24599 => "11001001",
                     24600 => "00000110",
                     24601 => "11010000",
                     24602 => "00000011",
                     24603 => "00100000",
                     24604 => "10010110",
                     24605 => "11100001",
                     24606 => "10101001",
                     24607 => "00000001",
                     24608 => "00100000",
                     24609 => "00010011",
                     24610 => "11011010",
                     24611 => "11001001",
                     24612 => "00001001",
                     24613 => "10010000",
                     24614 => "00010000",
                     24615 => "11001001",
                     24616 => "00010001",
                     24617 => "10110000",
                     24618 => "00001100",
                     24619 => "11001001",
                     24620 => "00001010",
                     24621 => "10010000",
                     24622 => "00000100",
                     24623 => "11001001",
                     24624 => "00001101",
                     24625 => "10010000",
                     24626 => "00000100",
                     24627 => "00101001",
                     24628 => "00000001",
                     24629 => "10010101",
                     24630 => "00010110",
                     24631 => "10110101",
                     24632 => "00011110",
                     24633 => "00101001",
                     24634 => "11110000",
                     24635 => "00001001",
                     24636 => "00000010",
                     24637 => "10010101",
                     24638 => "00011110",
                     24639 => "11010110",
                     24640 => "11001111",
                     24641 => "11010110",
                     24642 => "11001111",
                     24643 => "10110101",
                     24644 => "00010110",
                     24645 => "11001001",
                     24646 => "00000111",
                     24647 => "11110000",
                     24648 => "00000111",
                     24649 => "10101001",
                     24650 => "11111101",
                     24651 => "10101100",
                     24652 => "01001110",
                     24653 => "00000111",
                     24654 => "11010000",
                     24655 => "00000010",
                     24656 => "10101001",
                     24657 => "11111111",
                     24658 => "10010101",
                     24659 => "10100000",
                     24660 => "10100000",
                     24661 => "00000001",
                     24662 => "00100000",
                     24663 => "01001011",
                     24664 => "11100001",
                     24665 => "00010000",
                     24666 => "00000001",
                     24667 => "11001000",
                     24668 => "10110101",
                     24669 => "00010110",
                     24670 => "11001001",
                     24671 => "00110011",
                     24672 => "11110000",
                     24673 => "00000110",
                     24674 => "11001001",
                     24675 => "00001000",
                     24676 => "11110000",
                     24677 => "00000010",
                     24678 => "10010100",
                     24679 => "01000110",
                     24680 => "10001000",
                     24681 => "10111001",
                     24682 => "11000111",
                     24683 => "11011111",
                     24684 => "10010101",
                     24685 => "01011000",
                     24686 => "01100000",
                     24687 => "10100101",
                     24688 => "00000100",
                     24689 => "00111000",
                     24690 => "11101001",
                     24691 => "00001000",
                     24692 => "11001001",
                     24693 => "00000101",
                     24694 => "10110000",
                     24695 => "01110010",
                     24696 => "10110101",
                     24697 => "00011110",
                     24698 => "00101001",
                     24699 => "01000000",
                     24700 => "11010000",
                     24701 => "01010111",
                     24702 => "10110101",
                     24703 => "00011110",
                     24704 => "00001010",
                     24705 => "10010000",
                     24706 => "00000011",
                     24707 => "01001100",
                     24708 => "00000110",
                     24709 => "11100001",
                     24710 => "10110101",
                     24711 => "00011110",
                     24712 => "11110000",
                     24713 => "11111001",
                     24714 => "11001001",
                     24715 => "00000101",
                     24716 => "11110000",
                     24717 => "00011111",
                     24718 => "11001001",
                     24719 => "00000011",
                     24720 => "10110000",
                     24721 => "00011010",
                     24722 => "10110101",
                     24723 => "00011110",
                     24724 => "11001001",
                     24725 => "00000010",
                     24726 => "11010000",
                     24727 => "00010101",
                     24728 => "10101001",
                     24729 => "00010000",
                     24730 => "10110100",
                     24731 => "00010110",
                     24732 => "11000000",
                     24733 => "00010010",
                     24734 => "11010000",
                     24735 => "00000010",
                     24736 => "10101001",
                     24737 => "00000000",
                     24738 => "10011101",
                     24739 => "10010110",
                     24740 => "00000111",
                     24741 => "10101001",
                     24742 => "00000011",
                     24743 => "10010101",
                     24744 => "00011110",
                     24745 => "00100000",
                     24746 => "01010111",
                     24747 => "11100001",
                     24748 => "01100000",
                     24749 => "10110101",
                     24750 => "00010110",
                     24751 => "11001001",
                     24752 => "00000110",
                     24753 => "11110000",
                     24754 => "00100010",
                     24755 => "11001001",
                     24756 => "00010010",
                     24757 => "11010000",
                     24758 => "00001110",
                     24759 => "10101001",
                     24760 => "00000001",
                     24761 => "10010101",
                     24762 => "01000110",
                     24763 => "10101001",
                     24764 => "00001000",
                     24765 => "10010101",
                     24766 => "01011000",
                     24767 => "10100101",
                     24768 => "00001001",
                     24769 => "00101001",
                     24770 => "00000111",
                     24771 => "11110000",
                     24772 => "00010000",
                     24773 => "10100000",
                     24774 => "00000001",
                     24775 => "00100000",
                     24776 => "01001011",
                     24777 => "11100001",
                     24778 => "00010000",
                     24779 => "00000001",
                     24780 => "11001000",
                     24781 => "10011000",
                     24782 => "11010101",
                     24783 => "01000110",
                     24784 => "11010000",
                     24785 => "00000011",
                     24786 => "00100000",
                     24787 => "00101100",
                     24788 => "11100001",
                     24789 => "00100000",
                     24790 => "01010111",
                     24791 => "11100001",
                     24792 => "10110101",
                     24793 => "00011110",
                     24794 => "00101001",
                     24795 => "10000000",
                     24796 => "11010000",
                     24797 => "00000101",
                     24798 => "10101001",
                     24799 => "00000000",
                     24800 => "10010101",
                     24801 => "00011110",
                     24802 => "01100000",
                     24803 => "10110101",
                     24804 => "00011110",
                     24805 => "00101001",
                     24806 => "10111111",
                     24807 => "10010101",
                     24808 => "00011110",
                     24809 => "01100000",
                     24810 => "10110101",
                     24811 => "00010110",
                     24812 => "11001001",
                     24813 => "00000011",
                     24814 => "11010000",
                     24815 => "00000100",
                     24816 => "10110101",
                     24817 => "00011110",
                     24818 => "11110000",
                     24819 => "00111000",
                     24820 => "10110101",
                     24821 => "00011110",
                     24822 => "10101000",
                     24823 => "00001010",
                     24824 => "10010000",
                     24825 => "00000111",
                     24826 => "10110101",
                     24827 => "00011110",
                     24828 => "00001001",
                     24829 => "01000000",
                     24830 => "01001100",
                     24831 => "00000100",
                     24832 => "11100001",
                     24833 => "10111001",
                     24834 => "11000001",
                     24835 => "11011111",
                     24836 => "10010101",
                     24837 => "00011110",
                     24838 => "10110101",
                     24839 => "11001111",
                     24840 => "11001001",
                     24841 => "00100000",
                     24842 => "10010000",
                     24843 => "00011111",
                     24844 => "10100000",
                     24845 => "00010110",
                     24846 => "10101001",
                     24847 => "00000010",
                     24848 => "10000101",
                     24849 => "11101011",
                     24850 => "10100101",
                     24851 => "11101011",
                     24852 => "11010101",
                     24853 => "01000110",
                     24854 => "11010000",
                     24855 => "00001100",
                     24856 => "10101001",
                     24857 => "00000001",
                     24858 => "00100000",
                     24859 => "10010000",
                     24860 => "11100011",
                     24861 => "11110000",
                     24862 => "00000101",
                     24863 => "00100000",
                     24864 => "10111101",
                     24865 => "11100001",
                     24866 => "11010000",
                     24867 => "00001000",
                     24868 => "11000110",
                     24869 => "11101011",
                     24870 => "11001000",
                     24871 => "11000000",
                     24872 => "00011000",
                     24873 => "10010000",
                     24874 => "11100111",
                     24875 => "01100000",
                     24876 => "11100000",
                     24877 => "00000101",
                     24878 => "11110000",
                     24879 => "00001001",
                     24880 => "10110101",
                     24881 => "00011110",
                     24882 => "00001010",
                     24883 => "10010000",
                     24884 => "00000100",
                     24885 => "10101001",
                     24886 => "00000010",
                     24887 => "10000101",
                     24888 => "11111111",
                     24889 => "10110101",
                     24890 => "00010110",
                     24891 => "11001001",
                     24892 => "00000101",
                     24893 => "11010000",
                     24894 => "00001001",
                     24895 => "10101001",
                     24896 => "00000000",
                     24897 => "10000101",
                     24898 => "00000000",
                     24899 => "10100000",
                     24900 => "11111010",
                     24901 => "01001100",
                     24902 => "00111101",
                     24903 => "11001010",
                     24904 => "01001100",
                     24905 => "00111000",
                     24906 => "11011011",
                     24907 => "10110101",
                     24908 => "10000111",
                     24909 => "00111000",
                     24910 => "11100101",
                     24911 => "10000110",
                     24912 => "10000101",
                     24913 => "00000000",
                     24914 => "10110101",
                     24915 => "01101110",
                     24916 => "11100101",
                     24917 => "01101101",
                     24918 => "01100000",
                     24919 => "00100000",
                     24920 => "01101001",
                     24921 => "11000011",
                     24922 => "10110101",
                     24923 => "11001111",
                     24924 => "00101001",
                     24925 => "11110000",
                     24926 => "00001001",
                     24927 => "00001000",
                     24928 => "10010101",
                     24929 => "11001111",
                     24930 => "01100000",
                     24931 => "10110101",
                     24932 => "11001111",
                     24933 => "00011000",
                     24934 => "01101001",
                     24935 => "00111110",
                     24936 => "11001001",
                     24937 => "01000100",
                     24938 => "01100000",
                     24939 => "00100000",
                     24940 => "01100011",
                     24941 => "11100001",
                     24942 => "10010000",
                     24943 => "00011010",
                     24944 => "10110101",
                     24945 => "10100000",
                     24946 => "00011000",
                     24947 => "01101001",
                     24948 => "00000010",
                     24949 => "11001001",
                     24950 => "00000011",
                     24951 => "10010000",
                     24952 => "00010001",
                     24953 => "00100000",
                     24954 => "10110110",
                     24955 => "11100001",
                     24956 => "11110000",
                     24957 => "00001100",
                     24958 => "00100000",
                     24959 => "10111101",
                     24960 => "11100001",
                     24961 => "11110000",
                     24962 => "00000111",
                     24963 => "00100000",
                     24964 => "01010111",
                     24965 => "11100001",
                     24966 => "10101001",
                     24967 => "11111101",
                     24968 => "10010101",
                     24969 => "10100000",
                     24970 => "01001100",
                     24971 => "00000110",
                     24972 => "11100001",
                     24973 => "00100000",
                     24974 => "10110110",
                     24975 => "11100001",
                     24976 => "11110000",
                     24977 => "00011101",
                     24978 => "11001001",
                     24979 => "00100011",
                     24980 => "11010000",
                     24981 => "00001000",
                     24982 => "00100000",
                     24983 => "10010101",
                     24984 => "11010111",
                     24985 => "10101001",
                     24986 => "11111100",
                     24987 => "10010101",
                     24988 => "10100000",
                     24989 => "01100000",
                     24990 => "10111101",
                     24991 => "10001010",
                     24992 => "00000111",
                     24993 => "11010000",
                     24994 => "00001100",
                     24995 => "10110101",
                     24996 => "00011110",
                     24997 => "00101001",
                     24998 => "10001000",
                     24999 => "10010101",
                     25000 => "00011110",
                     25001 => "00100000",
                     25002 => "01010111",
                     25003 => "11100001",
                     25004 => "01001100",
                     25005 => "00000110",
                     25006 => "11100001",
                     25007 => "10110101",
                     25008 => "00011110",
                     25009 => "00001001",
                     25010 => "00000001",
                     25011 => "10010101",
                     25012 => "00011110",
                     25013 => "01100000",
                     25014 => "10101001",
                     25015 => "00000000",
                     25016 => "10100000",
                     25017 => "00010101",
                     25018 => "01001100",
                     25019 => "10010000",
                     25020 => "11100011",
                     25021 => "11001001",
                     25022 => "00100110",
                     25023 => "11110000",
                     25024 => "00001110",
                     25025 => "11001001",
                     25026 => "11000010",
                     25027 => "11110000",
                     25028 => "00001010",
                     25029 => "11001001",
                     25030 => "11000011",
                     25031 => "11110000",
                     25032 => "00000110",
                     25033 => "11001001",
                     25034 => "01011111",
                     25035 => "11110000",
                     25036 => "00000010",
                     25037 => "11001001",
                     25038 => "01100000",
                     25039 => "01100000",
                     25040 => "10110101",
                     25041 => "11010101",
                     25042 => "11001001",
                     25043 => "00011000",
                     25044 => "10010000",
                     25045 => "00100001",
                     25046 => "00100000",
                     25047 => "10100100",
                     25048 => "11100011",
                     25049 => "11110000",
                     25050 => "00011100",
                     25051 => "00100000",
                     25052 => "10111101",
                     25053 => "11100001",
                     25054 => "11110000",
                     25055 => "00010111",
                     25056 => "10110101",
                     25057 => "10100110",
                     25058 => "00110000",
                     25059 => "00011000",
                     25060 => "10110101",
                     25061 => "00111010",
                     25062 => "11010000",
                     25063 => "00010100",
                     25064 => "10101001",
                     25065 => "11111101",
                     25066 => "10010101",
                     25067 => "10100110",
                     25068 => "10101001",
                     25069 => "00000001",
                     25070 => "10010101",
                     25071 => "00111010",
                     25072 => "10110101",
                     25073 => "11010101",
                     25074 => "00101001",
                     25075 => "11111000",
                     25076 => "10010101",
                     25077 => "11010101",
                     25078 => "01100000",
                     25079 => "10101001",
                     25080 => "00000000",
                     25081 => "10010101",
                     25082 => "00111010",
                     25083 => "01100000",
                     25084 => "10101001",
                     25085 => "10000000",
                     25086 => "10010101",
                     25087 => "00100100",
                     25088 => "10101001",
                     25089 => "00000010",
                     25090 => "10000101",
                     25091 => "11111111",
                     25092 => "01100000",
                     25093 => "00000010",
                     25094 => "00001000",
                     25095 => "00001110",
                     25096 => "00100000",
                     25097 => "00000011",
                     25098 => "00010100",
                     25099 => "00001101",
                     25100 => "00100000",
                     25101 => "00000010",
                     25102 => "00010100",
                     25103 => "00001110",
                     25104 => "00100000",
                     25105 => "00000010",
                     25106 => "00001001",
                     25107 => "00001110",
                     25108 => "00010101",
                     25109 => "00000000",
                     25110 => "00000000",
                     25111 => "00011000",
                     25112 => "00000110",
                     25113 => "00000000",
                     25114 => "00000000",
                     25115 => "00100000",
                     25116 => "00001101",
                     25117 => "00000000",
                     25118 => "00000000",
                     25119 => "00110000",
                     25120 => "00001101",
                     25121 => "00000000",
                     25122 => "00000000",
                     25123 => "00001000",
                     25124 => "00001000",
                     25125 => "00000110",
                     25126 => "00000100",
                     25127 => "00001010",
                     25128 => "00001000",
                     25129 => "00000011",
                     25130 => "00001100",
                     25131 => "00001101",
                     25132 => "00010100",
                     25133 => "00000000",
                     25134 => "00000010",
                     25135 => "00010000",
                     25136 => "00010101",
                     25137 => "00000100",
                     25138 => "00000100",
                     25139 => "00001100",
                     25140 => "00011100",
                     25141 => "10001010",
                     25142 => "00011000",
                     25143 => "01101001",
                     25144 => "00000111",
                     25145 => "10101010",
                     25146 => "10100000",
                     25147 => "00000010",
                     25148 => "11010000",
                     25149 => "00000111",
                     25150 => "10001010",
                     25151 => "00011000",
                     25152 => "01101001",
                     25153 => "00001001",
                     25154 => "10101010",
                     25155 => "10100000",
                     25156 => "00000110",
                     25157 => "00100000",
                     25158 => "10100100",
                     25159 => "11100010",
                     25160 => "01001100",
                     25161 => "11100110",
                     25162 => "11100010",
                     25163 => "10100000",
                     25164 => "01001000",
                     25165 => "10000100",
                     25166 => "00000000",
                     25167 => "10100000",
                     25168 => "01000100",
                     25169 => "01001100",
                     25170 => "01011010",
                     25171 => "11100010",
                     25172 => "10100000",
                     25173 => "00001000",
                     25174 => "10000100",
                     25175 => "00000000",
                     25176 => "10100000",
                     25177 => "00000100",
                     25178 => "10110101",
                     25179 => "10000111",
                     25180 => "00111000",
                     25181 => "11101101",
                     25182 => "00011100",
                     25183 => "00000111",
                     25184 => "10000101",
                     25185 => "00000001",
                     25186 => "10110101",
                     25187 => "01101110",
                     25188 => "11101101",
                     25189 => "00011010",
                     25190 => "00000111",
                     25191 => "00110000",
                     25192 => "00000110",
                     25193 => "00000101",
                     25194 => "00000001",
                     25195 => "11110000",
                     25196 => "00000010",
                     25197 => "10100100",
                     25198 => "00000000",
                     25199 => "10011000",
                     25200 => "00101101",
                     25201 => "11010001",
                     25202 => "00000011",
                     25203 => "10011101",
                     25204 => "11011000",
                     25205 => "00000011",
                     25206 => "11010000",
                     25207 => "00011001",
                     25208 => "01001100",
                     25209 => "10000100",
                     25210 => "11100010",
                     25211 => "11101000",
                     25212 => "00100000",
                     25213 => "11111101",
                     25214 => "11110001",
                     25215 => "11001010",
                     25216 => "11001001",
                     25217 => "11111110",
                     25218 => "10110000",
                     25219 => "00001101",
                     25220 => "10001010",
                     25221 => "00011000",
                     25222 => "01101001",
                     25223 => "00000001",
                     25224 => "10101010",
                     25225 => "10100000",
                     25226 => "00000001",
                     25227 => "00100000",
                     25228 => "10100100",
                     25229 => "11100010",
                     25230 => "01001100",
                     25231 => "11100110",
                     25232 => "11100010",
                     25233 => "10001010",
                     25234 => "00001010",
                     25235 => "00001010",
                     25236 => "10101000",
                     25237 => "10101001",
                     25238 => "11111111",
                     25239 => "10011001",
                     25240 => "10110000",
                     25241 => "00000100",
                     25242 => "10011001",
                     25243 => "10110001",
                     25244 => "00000100",
                     25245 => "10011001",
                     25246 => "10110010",
                     25247 => "00000100",
                     25248 => "10011001",
                     25249 => "10110011",
                     25250 => "00000100",
                     25251 => "01100000",
                     25252 => "10000110",
                     25253 => "00000000",
                     25254 => "10111001",
                     25255 => "10111000",
                     25256 => "00000011",
                     25257 => "10000101",
                     25258 => "00000010",
                     25259 => "10111001",
                     25260 => "10101101",
                     25261 => "00000011",
                     25262 => "10000101",
                     25263 => "00000001",
                     25264 => "10001010",
                     25265 => "00001010",
                     25266 => "00001010",
                     25267 => "01001000",
                     25268 => "10101000",
                     25269 => "10111101",
                     25270 => "10011001",
                     25271 => "00000100",
                     25272 => "00001010",
                     25273 => "00001010",
                     25274 => "10101010",
                     25275 => "10100101",
                     25276 => "00000001",
                     25277 => "00011000",
                     25278 => "01111101",
                     25279 => "00000101",
                     25280 => "11100010",
                     25281 => "10011001",
                     25282 => "10101100",
                     25283 => "00000100",
                     25284 => "10100101",
                     25285 => "00000001",
                     25286 => "00011000",
                     25287 => "01111101",
                     25288 => "00000111",
                     25289 => "11100010",
                     25290 => "10011001",
                     25291 => "10101110",
                     25292 => "00000100",
                     25293 => "11101000",
                     25294 => "11001000",
                     25295 => "10100101",
                     25296 => "00000010",
                     25297 => "00011000",
                     25298 => "01111101",
                     25299 => "00000101",
                     25300 => "11100010",
                     25301 => "10011001",
                     25302 => "10101100",
                     25303 => "00000100",
                     25304 => "10100101",
                     25305 => "00000010",
                     25306 => "00011000",
                     25307 => "01111101",
                     25308 => "00000111",
                     25309 => "11100010",
                     25310 => "10011001",
                     25311 => "10101110",
                     25312 => "00000100",
                     25313 => "01101000",
                     25314 => "10101000",
                     25315 => "10100110",
                     25316 => "00000000",
                     25317 => "01100000",
                     25318 => "10101101",
                     25319 => "00011100",
                     25320 => "00000111",
                     25321 => "00011000",
                     25322 => "01101001",
                     25323 => "10000000",
                     25324 => "10000101",
                     25325 => "00000010",
                     25326 => "10101101",
                     25327 => "00011010",
                     25328 => "00000111",
                     25329 => "01101001",
                     25330 => "00000000",
                     25331 => "10000101",
                     25332 => "00000001",
                     25333 => "10110101",
                     25334 => "10000110",
                     25335 => "11000101",
                     25336 => "00000010",
                     25337 => "10110101",
                     25338 => "01101101",
                     25339 => "11100101",
                     25340 => "00000001",
                     25341 => "10010000",
                     25342 => "00010101",
                     25343 => "10111001",
                     25344 => "10101110",
                     25345 => "00000100",
                     25346 => "00110000",
                     25347 => "00001101",
                     25348 => "10101001",
                     25349 => "11111111",
                     25350 => "10111110",
                     25351 => "10101100",
                     25352 => "00000100",
                     25353 => "00110000",
                     25354 => "00000011",
                     25355 => "10011001",
                     25356 => "10101100",
                     25357 => "00000100",
                     25358 => "10011001",
                     25359 => "10101110",
                     25360 => "00000100",
                     25361 => "10100110",
                     25362 => "00001000",
                     25363 => "01100000",
                     25364 => "10111001",
                     25365 => "10101100",
                     25366 => "00000100",
                     25367 => "00010000",
                     25368 => "00010001",
                     25369 => "11001001",
                     25370 => "10100000",
                     25371 => "10010000",
                     25372 => "00001101",
                     25373 => "10101001",
                     25374 => "00000000",
                     25375 => "10111110",
                     25376 => "10101110",
                     25377 => "00000100",
                     25378 => "00010000",
                     25379 => "00000011",
                     25380 => "10011001",
                     25381 => "10101110",
                     25382 => "00000100",
                     25383 => "10011001",
                     25384 => "10101100",
                     25385 => "00000100",
                     25386 => "10100110",
                     25387 => "00001000",
                     25388 => "01100000",
                     25389 => "10100010",
                     25390 => "00000000",
                     25391 => "10000100",
                     25392 => "00000110",
                     25393 => "10101001",
                     25394 => "00000001",
                     25395 => "10000101",
                     25396 => "00000111",
                     25397 => "10111001",
                     25398 => "10101100",
                     25399 => "00000100",
                     25400 => "11011101",
                     25401 => "10101100",
                     25402 => "00000100",
                     25403 => "10110000",
                     25404 => "00101010",
                     25405 => "11011101",
                     25406 => "10101110",
                     25407 => "00000100",
                     25408 => "10010000",
                     25409 => "00010010",
                     25410 => "11110000",
                     25411 => "01000010",
                     25412 => "10111001",
                     25413 => "10101110",
                     25414 => "00000100",
                     25415 => "11011001",
                     25416 => "10101100",
                     25417 => "00000100",
                     25418 => "10010000",
                     25419 => "00111010",
                     25420 => "11011101",
                     25421 => "10101100",
                     25422 => "00000100",
                     25423 => "10110000",
                     25424 => "00110101",
                     25425 => "10100100",
                     25426 => "00000110",
                     25427 => "01100000",
                     25428 => "10111101",
                     25429 => "10101110",
                     25430 => "00000100",
                     25431 => "11011101",
                     25432 => "10101100",
                     25433 => "00000100",
                     25434 => "10010000",
                     25435 => "00101010",
                     25436 => "10111001",
                     25437 => "10101110",
                     25438 => "00000100",
                     25439 => "11011101",
                     25440 => "10101100",
                     25441 => "00000100",
                     25442 => "10110000",
                     25443 => "00100010",
                     25444 => "10100100",
                     25445 => "00000110",
                     25446 => "01100000",
                     25447 => "11011101",
                     25448 => "10101100",
                     25449 => "00000100",
                     25450 => "11110000",
                     25451 => "00011010",
                     25452 => "11011101",
                     25453 => "10101110",
                     25454 => "00000100",
                     25455 => "10010000",
                     25456 => "00010101",
                     25457 => "11110000",
                     25458 => "00010011",
                     25459 => "11011001",
                     25460 => "10101110",
                     25461 => "00000100",
                     25462 => "10010000",
                     25463 => "00001010",
                     25464 => "11110000",
                     25465 => "00001000",
                     25466 => "10111001",
                     25467 => "10101110",
                     25468 => "00000100",
                     25469 => "11011101",
                     25470 => "10101100",
                     25471 => "00000100",
                     25472 => "10110000",
                     25473 => "00000100",
                     25474 => "00011000",
                     25475 => "10100100",
                     25476 => "00000110",
                     25477 => "01100000",
                     25478 => "11101000",
                     25479 => "11001000",
                     25480 => "11000110",
                     25481 => "00000111",
                     25482 => "00010000",
                     25483 => "10101001",
                     25484 => "00111000",
                     25485 => "10100100",
                     25486 => "00000110",
                     25487 => "01100000",
                     25488 => "01001000",
                     25489 => "10001010",
                     25490 => "00011000",
                     25491 => "01101001",
                     25492 => "00000001",
                     25493 => "10101010",
                     25494 => "01101000",
                     25495 => "01001100",
                     25496 => "10101101",
                     25497 => "11100011",
                     25498 => "10001010",
                     25499 => "00011000",
                     25500 => "01101001",
                     25501 => "00001101",
                     25502 => "10101010",
                     25503 => "10100000",
                     25504 => "00011011",
                     25505 => "01001100",
                     25506 => "10101011",
                     25507 => "11100011",
                     25508 => "10100000",
                     25509 => "00011010",
                     25510 => "10001010",
                     25511 => "00011000",
                     25512 => "01101001",
                     25513 => "00000111",
                     25514 => "10101010",
                     25515 => "10101001",
                     25516 => "00000000",
                     25517 => "00100000",
                     25518 => "11111000",
                     25519 => "11100011",
                     25520 => "10100110",
                     25521 => "00001000",
                     25522 => "11001001",
                     25523 => "00000000",
                     25524 => "01100000",
                     25525 => "00000000",
                     25526 => "00000111",
                     25527 => "00001110",
                     25528 => "00001000",
                     25529 => "00000011",
                     25530 => "00001100",
                     25531 => "00000010",
                     25532 => "00000010",
                     25533 => "00001101",
                     25534 => "00001101",
                     25535 => "00001000",
                     25536 => "00000011",
                     25537 => "00001100",
                     25538 => "00000010",
                     25539 => "00000010",
                     25540 => "00001101",
                     25541 => "00001101",
                     25542 => "00001000",
                     25543 => "00000011",
                     25544 => "00001100",
                     25545 => "00000010",
                     25546 => "00000010",
                     25547 => "00001101",
                     25548 => "00001101",
                     25549 => "00001000",
                     25550 => "00000000",
                     25551 => "00010000",
                     25552 => "00000100",
                     25553 => "00010100",
                     25554 => "00000100",
                     25555 => "00000100",
                     25556 => "00000100",
                     25557 => "00100000",
                     25558 => "00100000",
                     25559 => "00001000",
                     25560 => "00011000",
                     25561 => "00001000",
                     25562 => "00011000",
                     25563 => "00000010",
                     25564 => "00100000",
                     25565 => "00100000",
                     25566 => "00001000",
                     25567 => "00011000",
                     25568 => "00001000",
                     25569 => "00011000",
                     25570 => "00010010",
                     25571 => "00100000",
                     25572 => "00100000",
                     25573 => "00011000",
                     25574 => "00011000",
                     25575 => "00011000",
                     25576 => "00011000",
                     25577 => "00011000",
                     25578 => "00010100",
                     25579 => "00010100",
                     25580 => "00000110",
                     25581 => "00000110",
                     25582 => "00001000",
                     25583 => "00010000",
                     25584 => "11001000",
                     25585 => "10101001",
                     25586 => "00000000",
                     25587 => "00101100",
                     25588 => "10101001",
                     25589 => "00000001",
                     25590 => "10100010",
                     25591 => "00000000",
                     25592 => "01001000",
                     25593 => "10000100",
                     25594 => "00000100",
                     25595 => "10111001",
                     25596 => "10111000",
                     25597 => "11100011",
                     25598 => "00011000",
                     25599 => "01110101",
                     25600 => "10000110",
                     25601 => "10000101",
                     25602 => "00000101",
                     25603 => "10110101",
                     25604 => "01101101",
                     25605 => "01101001",
                     25606 => "00000000",
                     25607 => "00101001",
                     25608 => "00000001",
                     25609 => "01001010",
                     25610 => "00000101",
                     25611 => "00000101",
                     25612 => "01101010",
                     25613 => "01001010",
                     25614 => "01001010",
                     25615 => "01001010",
                     25616 => "00100000",
                     25617 => "11100011",
                     25618 => "10011011",
                     25619 => "10100100",
                     25620 => "00000100",
                     25621 => "10110101",
                     25622 => "11001110",
                     25623 => "00011000",
                     25624 => "01111001",
                     25625 => "11010100",
                     25626 => "11100011",
                     25627 => "00101001",
                     25628 => "11110000",
                     25629 => "00111000",
                     25630 => "11101001",
                     25631 => "00100000",
                     25632 => "10000101",
                     25633 => "00000010",
                     25634 => "10101000",
                     25635 => "10110001",
                     25636 => "00000110",
                     25637 => "10000101",
                     25638 => "00000011",
                     25639 => "10100100",
                     25640 => "00000100",
                     25641 => "01101000",
                     25642 => "11010000",
                     25643 => "00000101",
                     25644 => "10110101",
                     25645 => "11001110",
                     25646 => "01001100",
                     25647 => "00110011",
                     25648 => "11100100",
                     25649 => "10110101",
                     25650 => "10000110",
                     25651 => "00101001",
                     25652 => "00001111",
                     25653 => "10000101",
                     25654 => "00000100",
                     25655 => "10100101",
                     25656 => "00000011",
                     25657 => "01100000",
                     25658 => "00000000",
                     25659 => "00110000",
                     25660 => "10000100",
                     25661 => "00000000",
                     25662 => "10101101",
                     25663 => "10111001",
                     25664 => "00000011",
                     25665 => "00011000",
                     25666 => "01111001",
                     25667 => "00111010",
                     25668 => "11100100",
                     25669 => "10111110",
                     25670 => "10011010",
                     25671 => "00000011",
                     25672 => "10111100",
                     25673 => "11100101",
                     25674 => "00000110",
                     25675 => "10000100",
                     25676 => "00000010",
                     25677 => "00100000",
                     25678 => "10110101",
                     25679 => "11100100",
                     25680 => "10101101",
                     25681 => "10101110",
                     25682 => "00000011",
                     25683 => "10011001",
                     25684 => "00000011",
                     25685 => "00000010",
                     25686 => "10011001",
                     25687 => "00001011",
                     25688 => "00000010",
                     25689 => "10011001",
                     25690 => "00010011",
                     25691 => "00000010",
                     25692 => "00011000",
                     25693 => "01101001",
                     25694 => "00000110",
                     25695 => "10011001",
                     25696 => "00000111",
                     25697 => "00000010",
                     25698 => "10011001",
                     25699 => "00001111",
                     25700 => "00000010",
                     25701 => "10011001",
                     25702 => "00010111",
                     25703 => "00000010",
                     25704 => "10101001",
                     25705 => "00100001",
                     25706 => "10011001",
                     25707 => "00000010",
                     25708 => "00000010",
                     25709 => "10011001",
                     25710 => "00001010",
                     25711 => "00000010",
                     25712 => "10011001",
                     25713 => "00010010",
                     25714 => "00000010",
                     25715 => "00001001",
                     25716 => "01000000",
                     25717 => "10011001",
                     25718 => "00000110",
                     25719 => "00000010",
                     25720 => "10011001",
                     25721 => "00001110",
                     25722 => "00000010",
                     25723 => "10011001",
                     25724 => "00010110",
                     25725 => "00000010",
                     25726 => "10100010",
                     25727 => "00000101",
                     25728 => "10101001",
                     25729 => "11100001",
                     25730 => "10011001",
                     25731 => "00000001",
                     25732 => "00000010",
                     25733 => "11001000",
                     25734 => "11001000",
                     25735 => "11001000",
                     25736 => "11001000",
                     25737 => "11001010",
                     25738 => "00010000",
                     25739 => "11110100",
                     25740 => "10100100",
                     25741 => "00000010",
                     25742 => "10100101",
                     25743 => "00000000",
                     25744 => "11010000",
                     25745 => "00000101",
                     25746 => "10101001",
                     25747 => "11100000",
                     25748 => "10011001",
                     25749 => "00000001",
                     25750 => "00000010",
                     25751 => "10100010",
                     25752 => "00000000",
                     25753 => "10101101",
                     25754 => "10011101",
                     25755 => "00000011",
                     25756 => "00111000",
                     25757 => "11111001",
                     25758 => "00000000",
                     25759 => "00000010",
                     25760 => "11001001",
                     25761 => "01100100",
                     25762 => "10010000",
                     25763 => "00000101",
                     25764 => "10101001",
                     25765 => "11111000",
                     25766 => "10011001",
                     25767 => "00000000",
                     25768 => "00000010",
                     25769 => "11001000",
                     25770 => "11001000",
                     25771 => "11001000",
                     25772 => "11001000",
                     25773 => "11101000",
                     25774 => "11100000",
                     25775 => "00000110",
                     25776 => "11010000",
                     25777 => "11100111",
                     25778 => "10100100",
                     25779 => "00000000",
                     25780 => "01100000",
                     25781 => "10100010",
                     25782 => "00000110",
                     25783 => "10011001",
                     25784 => "00000000",
                     25785 => "00000010",
                     25786 => "00011000",
                     25787 => "01101001",
                     25788 => "00001000",
                     25789 => "11001000",
                     25790 => "11001000",
                     25791 => "11001000",
                     25792 => "11001000",
                     25793 => "11001010",
                     25794 => "11010000",
                     25795 => "11110011",
                     25796 => "10100100",
                     25797 => "00000010",
                     25798 => "01100000",
                     25799 => "00000100",
                     25800 => "00000000",
                     25801 => "00000100",
                     25802 => "00000000",
                     25803 => "00000000",
                     25804 => "00000100",
                     25805 => "00000000",
                     25806 => "00000100",
                     25807 => "00000000",
                     25808 => "00001000",
                     25809 => "00000000",
                     25810 => "00001000",
                     25811 => "00001000",
                     25812 => "00000000",
                     25813 => "00001000",
                     25814 => "00000000",
                     25815 => "10000000",
                     25816 => "10000010",
                     25817 => "10000001",
                     25818 => "10000011",
                     25819 => "10000001",
                     25820 => "10000011",
                     25821 => "10000000",
                     25822 => "10000010",
                     25823 => "00000011",
                     25824 => "00000011",
                     25825 => "11000011",
                     25826 => "11000011",
                     25827 => "10111100",
                     25828 => "11110011",
                     25829 => "00000110",
                     25830 => "10101101",
                     25831 => "01000111",
                     25832 => "00000111",
                     25833 => "11010000",
                     25834 => "00001000",
                     25835 => "10110101",
                     25836 => "00101010",
                     25837 => "00101001",
                     25838 => "01111111",
                     25839 => "11001001",
                     25840 => "00000001",
                     25841 => "11110000",
                     25842 => "00000100",
                     25843 => "10100010",
                     25844 => "00000000",
                     25845 => "11110000",
                     25846 => "00000111",
                     25847 => "10100101",
                     25848 => "00001001",
                     25849 => "01001010",
                     25850 => "01001010",
                     25851 => "00101001",
                     25852 => "00000011",
                     25853 => "10101010",
                     25854 => "10101101",
                     25855 => "10111110",
                     25856 => "00000011",
                     25857 => "00011000",
                     25858 => "01111101",
                     25859 => "11001011",
                     25860 => "11100100",
                     25861 => "10011001",
                     25862 => "00000000",
                     25863 => "00000010",
                     25864 => "00011000",
                     25865 => "01111101",
                     25866 => "11010011",
                     25867 => "11100100",
                     25868 => "10011001",
                     25869 => "00000100",
                     25870 => "00000010",
                     25871 => "10101101",
                     25872 => "10110011",
                     25873 => "00000011",
                     25874 => "00011000",
                     25875 => "01111101",
                     25876 => "11000111",
                     25877 => "11100100",
                     25878 => "10011001",
                     25879 => "00000011",
                     25880 => "00000010",
                     25881 => "00011000",
                     25882 => "01111101",
                     25883 => "11001111",
                     25884 => "11100100",
                     25885 => "10011001",
                     25886 => "00000111",
                     25887 => "00000010",
                     25888 => "10111101",
                     25889 => "11010111",
                     25890 => "11100100",
                     25891 => "10011001",
                     25892 => "00000001",
                     25893 => "00000010",
                     25894 => "10111101",
                     25895 => "11011011",
                     25896 => "11100100",
                     25897 => "10011001",
                     25898 => "00000101",
                     25899 => "00000010",
                     25900 => "10111101",
                     25901 => "11011111",
                     25902 => "11100100",
                     25903 => "10011001",
                     25904 => "00000010",
                     25905 => "00000010",
                     25906 => "10011001",
                     25907 => "00000110",
                     25908 => "00000010",
                     25909 => "10100110",
                     25910 => "00001000",
                     25911 => "10101101",
                     25912 => "11010110",
                     25913 => "00000011",
                     25914 => "00101001",
                     25915 => "11111100",
                     25916 => "11110000",
                     25917 => "00001001",
                     25918 => "10101001",
                     25919 => "00000000",
                     25920 => "10010101",
                     25921 => "00101010",
                     25922 => "10101001",
                     25923 => "11111000",
                     25924 => "00100000",
                     25925 => "11001000",
                     25926 => "11100101",
                     25927 => "01100000",
                     25928 => "11111001",
                     25929 => "01010000",
                     25930 => "11110111",
                     25931 => "01010000",
                     25932 => "11111010",
                     25933 => "11111011",
                     25934 => "11111000",
                     25935 => "11111011",
                     25936 => "11110110",
                     25937 => "11111011",
                     25938 => "10111100",
                     25939 => "11100101",
                     25940 => "00000110",
                     25941 => "10101101",
                     25942 => "10101110",
                     25943 => "00000011",
                     25944 => "10011001",
                     25945 => "00000011",
                     25946 => "00000010",
                     25947 => "00011000",
                     25948 => "01101001",
                     25949 => "00001000",
                     25950 => "10011001",
                     25951 => "00000111",
                     25952 => "00000010",
                     25953 => "10011001",
                     25954 => "00001011",
                     25955 => "00000010",
                     25956 => "00011000",
                     25957 => "01101001",
                     25958 => "00001100",
                     25959 => "10000101",
                     25960 => "00000101",
                     25961 => "10110101",
                     25962 => "11001111",
                     25963 => "00100000",
                     25964 => "11001000",
                     25965 => "11100101",
                     25966 => "01101001",
                     25967 => "00001000",
                     25968 => "10011001",
                     25969 => "00001000",
                     25970 => "00000010",
                     25971 => "10101101",
                     25972 => "00001101",
                     25973 => "00000001",
                     25974 => "10000101",
                     25975 => "00000010",
                     25976 => "10101001",
                     25977 => "00000001",
                     25978 => "10000101",
                     25979 => "00000011",
                     25980 => "10000101",
                     25981 => "00000100",
                     25982 => "10011001",
                     25983 => "00000010",
                     25984 => "00000010",
                     25985 => "10011001",
                     25986 => "00000110",
                     25987 => "00000010",
                     25988 => "10011001",
                     25989 => "00001010",
                     25990 => "00000010",
                     25991 => "10101001",
                     25992 => "01111110",
                     25993 => "10011001",
                     25994 => "00000001",
                     25995 => "00000010",
                     25996 => "10011001",
                     25997 => "00001001",
                     25998 => "00000010",
                     25999 => "10101001",
                     26000 => "01111111",
                     26001 => "10011001",
                     26002 => "00000101",
                     26003 => "00000010",
                     26004 => "10101101",
                     26005 => "00001111",
                     26006 => "00000111",
                     26007 => "11110000",
                     26008 => "00010101",
                     26009 => "10011000",
                     26010 => "00011000",
                     26011 => "01101001",
                     26012 => "00001100",
                     26013 => "10101000",
                     26014 => "10101101",
                     26015 => "00001111",
                     26016 => "00000001",
                     26017 => "00001010",
                     26018 => "10101010",
                     26019 => "10111101",
                     26020 => "01001000",
                     26021 => "11100101",
                     26022 => "10000101",
                     26023 => "00000000",
                     26024 => "10111101",
                     26025 => "01001001",
                     26026 => "11100101",
                     26027 => "00100000",
                     26028 => "10111001",
                     26029 => "11101011",
                     26030 => "10100110",
                     26031 => "00001000",
                     26032 => "10111100",
                     26033 => "11100101",
                     26034 => "00000110",
                     26035 => "10101101",
                     26036 => "11010001",
                     26037 => "00000011",
                     26038 => "00101001",
                     26039 => "00001110",
                     26040 => "11110000",
                     26041 => "00010100",
                     26042 => "10101001",
                     26043 => "11111000",
                     26044 => "10011001",
                     26045 => "00010100",
                     26046 => "00000010",
                     26047 => "10011001",
                     26048 => "00010000",
                     26049 => "00000010",
                     26050 => "10011001",
                     26051 => "00001100",
                     26052 => "00000010",
                     26053 => "10011001",
                     26054 => "00001000",
                     26055 => "00000010",
                     26056 => "10011001",
                     26057 => "00000100",
                     26058 => "00000010",
                     26059 => "10011001",
                     26060 => "00000000",
                     26061 => "00000010",
                     26062 => "01100000",
                     26063 => "10111100",
                     26064 => "11100101",
                     26065 => "00000110",
                     26066 => "10000100",
                     26067 => "00000010",
                     26068 => "11001000",
                     26069 => "11001000",
                     26070 => "11001000",
                     26071 => "10101101",
                     26072 => "10101110",
                     26073 => "00000011",
                     26074 => "00100000",
                     26075 => "10110101",
                     26076 => "11100100",
                     26077 => "10100110",
                     26078 => "00001000",
                     26079 => "10110101",
                     26080 => "11001111",
                     26081 => "00100000",
                     26082 => "11000010",
                     26083 => "11100101",
                     26084 => "10101100",
                     26085 => "01001110",
                     26086 => "00000111",
                     26087 => "11000000",
                     26088 => "00000011",
                     26089 => "11110000",
                     26090 => "00000101",
                     26091 => "10101100",
                     26092 => "11001100",
                     26093 => "00000110",
                     26094 => "11110000",
                     26095 => "00000010",
                     26096 => "10101001",
                     26097 => "11111000",
                     26098 => "10111100",
                     26099 => "11100101",
                     26100 => "00000110",
                     26101 => "10011001",
                     26102 => "00010000",
                     26103 => "00000010",
                     26104 => "10011001",
                     26105 => "00010100",
                     26106 => "00000010",
                     26107 => "10101001",
                     26108 => "01011011",
                     26109 => "10101110",
                     26110 => "01000011",
                     26111 => "00000111",
                     26112 => "11110000",
                     26113 => "00000010",
                     26114 => "10101001",
                     26115 => "01110101",
                     26116 => "10100110",
                     26117 => "00001000",
                     26118 => "11001000",
                     26119 => "00100000",
                     26120 => "10111100",
                     26121 => "11100101",
                     26122 => "10101001",
                     26123 => "00000010",
                     26124 => "11001000",
                     26125 => "00100000",
                     26126 => "10111100",
                     26127 => "11100101",
                     26128 => "11101000",
                     26129 => "00100000",
                     26130 => "11111101",
                     26131 => "11110001",
                     26132 => "11001010",
                     26133 => "10111100",
                     26134 => "11100101",
                     26135 => "00000110",
                     26136 => "00001010",
                     26137 => "01001000",
                     26138 => "10010000",
                     26139 => "00000101",
                     26140 => "10101001",
                     26141 => "11111000",
                     26142 => "10011001",
                     26143 => "00000000",
                     26144 => "00000010",
                     26145 => "01101000",
                     26146 => "00001010",
                     26147 => "01001000",
                     26148 => "10010000",
                     26149 => "00000101",
                     26150 => "10101001",
                     26151 => "11111000",
                     26152 => "10011001",
                     26153 => "00000100",
                     26154 => "00000010",
                     26155 => "01101000",
                     26156 => "00001010",
                     26157 => "01001000",
                     26158 => "10010000",
                     26159 => "00000101",
                     26160 => "10101001",
                     26161 => "11111000",
                     26162 => "10011001",
                     26163 => "00001000",
                     26164 => "00000010",
                     26165 => "01101000",
                     26166 => "00001010",
                     26167 => "01001000",
                     26168 => "10010000",
                     26169 => "00000101",
                     26170 => "10101001",
                     26171 => "11111000",
                     26172 => "10011001",
                     26173 => "00001100",
                     26174 => "00000010",
                     26175 => "01101000",
                     26176 => "00001010",
                     26177 => "01001000",
                     26178 => "10010000",
                     26179 => "00000101",
                     26180 => "10101001",
                     26181 => "11111000",
                     26182 => "10011001",
                     26183 => "00010000",
                     26184 => "00000010",
                     26185 => "01101000",
                     26186 => "00001010",
                     26187 => "10010000",
                     26188 => "00000101",
                     26189 => "10101001",
                     26190 => "11111000",
                     26191 => "10011001",
                     26192 => "00010100",
                     26193 => "00000010",
                     26194 => "10101101",
                     26195 => "11010001",
                     26196 => "00000011",
                     26197 => "00001010",
                     26198 => "10010000",
                     26199 => "00000011",
                     26200 => "00100000",
                     26201 => "10111010",
                     26202 => "11100101",
                     26203 => "01100000",
                     26204 => "10100101",
                     26205 => "00001001",
                     26206 => "01001010",
                     26207 => "10110000",
                     26208 => "00000010",
                     26209 => "11010110",
                     26210 => "11011011",
                     26211 => "10110101",
                     26212 => "11011011",
                     26213 => "00100000",
                     26214 => "11001000",
                     26215 => "11100101",
                     26216 => "10101101",
                     26217 => "10110011",
                     26218 => "00000011",
                     26219 => "10011001",
                     26220 => "00000011",
                     26221 => "00000010",
                     26222 => "00011000",
                     26223 => "01101001",
                     26224 => "00001000",
                     26225 => "10011001",
                     26226 => "00000111",
                     26227 => "00000010",
                     26228 => "10101001",
                     26229 => "00000010",
                     26230 => "10011001",
                     26231 => "00000010",
                     26232 => "00000010",
                     26233 => "10011001",
                     26234 => "00000110",
                     26235 => "00000010",
                     26236 => "10101001",
                     26237 => "11110111",
                     26238 => "10011001",
                     26239 => "00000001",
                     26240 => "00000010",
                     26241 => "10101001",
                     26242 => "11111011",
                     26243 => "10011001",
                     26244 => "00000101",
                     26245 => "00000010",
                     26246 => "01001100",
                     26247 => "11000100",
                     26248 => "11100110",
                     26249 => "01100000",
                     26250 => "01100001",
                     26251 => "01100010",
                     26252 => "01100011",
                     26253 => "10111100",
                     26254 => "11110011",
                     26255 => "00000110",
                     26256 => "10110101",
                     26257 => "00101010",
                     26258 => "11001001",
                     26259 => "00000010",
                     26260 => "10110000",
                     26261 => "11000110",
                     26262 => "10110101",
                     26263 => "11011011",
                     26264 => "10011001",
                     26265 => "00000000",
                     26266 => "00000010",
                     26267 => "00011000",
                     26268 => "01101001",
                     26269 => "00001000",
                     26270 => "10011001",
                     26271 => "00000100",
                     26272 => "00000010",
                     26273 => "10101101",
                     26274 => "10110011",
                     26275 => "00000011",
                     26276 => "10011001",
                     26277 => "00000011",
                     26278 => "00000010",
                     26279 => "10011001",
                     26280 => "00000111",
                     26281 => "00000010",
                     26282 => "10100101",
                     26283 => "00001001",
                     26284 => "01001010",
                     26285 => "00101001",
                     26286 => "00000011",
                     26287 => "10101010",
                     26288 => "10111101",
                     26289 => "10001001",
                     26290 => "11100110",
                     26291 => "11001000",
                     26292 => "00100000",
                     26293 => "11001000",
                     26294 => "11100101",
                     26295 => "10001000",
                     26296 => "10101001",
                     26297 => "00000010",
                     26298 => "10011001",
                     26299 => "00000010",
                     26300 => "00000010",
                     26301 => "10101001",
                     26302 => "10000010",
                     26303 => "10011001",
                     26304 => "00000110",
                     26305 => "00000010",
                     26306 => "10100110",
                     26307 => "00001000",
                     26308 => "01100000",
                     26309 => "01110110",
                     26310 => "01110111",
                     26311 => "01111000",
                     26312 => "01111001",
                     26313 => "11010110",
                     26314 => "11010110",
                     26315 => "11011001",
                     26316 => "11011001",
                     26317 => "10001101",
                     26318 => "10001101",
                     26319 => "11100100",
                     26320 => "11100100",
                     26321 => "01110110",
                     26322 => "01110111",
                     26323 => "01111000",
                     26324 => "01111001",
                     26325 => "00000010",
                     26326 => "00000001",
                     26327 => "00000010",
                     26328 => "00000001",
                     26329 => "10101100",
                     26330 => "11101010",
                     26331 => "00000110",
                     26332 => "10101101",
                     26333 => "10111001",
                     26334 => "00000011",
                     26335 => "00011000",
                     26336 => "01101001",
                     26337 => "00001000",
                     26338 => "10000101",
                     26339 => "00000010",
                     26340 => "10101101",
                     26341 => "10101110",
                     26342 => "00000011",
                     26343 => "10000101",
                     26344 => "00000101",
                     26345 => "10100110",
                     26346 => "00111001",
                     26347 => "10111101",
                     26348 => "11010101",
                     26349 => "11100110",
                     26350 => "00001101",
                     26351 => "11001010",
                     26352 => "00000011",
                     26353 => "10000101",
                     26354 => "00000100",
                     26355 => "10001010",
                     26356 => "01001000",
                     26357 => "00001010",
                     26358 => "00001010",
                     26359 => "10101010",
                     26360 => "10101001",
                     26361 => "00000001",
                     26362 => "10000101",
                     26363 => "00000111",
                     26364 => "10000101",
                     26365 => "00000011",
                     26366 => "10111101",
                     26367 => "11000101",
                     26368 => "11100110",
                     26369 => "10000101",
                     26370 => "00000000",
                     26371 => "10111101",
                     26372 => "11000110",
                     26373 => "11100110",
                     26374 => "00100000",
                     26375 => "10111001",
                     26376 => "11101011",
                     26377 => "11000110",
                     26378 => "00000111",
                     26379 => "00010000",
                     26380 => "11110001",
                     26381 => "10101100",
                     26382 => "11101010",
                     26383 => "00000110",
                     26384 => "01101000",
                     26385 => "11110000",
                     26386 => "00101111",
                     26387 => "11001001",
                     26388 => "00000011",
                     26389 => "11110000",
                     26390 => "00101011",
                     26391 => "10000101",
                     26392 => "00000000",
                     26393 => "10100101",
                     26394 => "00001001",
                     26395 => "01001010",
                     26396 => "00101001",
                     26397 => "00000011",
                     26398 => "00001101",
                     26399 => "11001010",
                     26400 => "00000011",
                     26401 => "10011001",
                     26402 => "00000010",
                     26403 => "00000010",
                     26404 => "10011001",
                     26405 => "00000110",
                     26406 => "00000010",
                     26407 => "10100110",
                     26408 => "00000000",
                     26409 => "11001010",
                     26410 => "11110000",
                     26411 => "00000110",
                     26412 => "10011001",
                     26413 => "00001010",
                     26414 => "00000010",
                     26415 => "10011001",
                     26416 => "00001110",
                     26417 => "00000010",
                     26418 => "10111001",
                     26419 => "00000110",
                     26420 => "00000010",
                     26421 => "00001001",
                     26422 => "01000000",
                     26423 => "10011001",
                     26424 => "00000110",
                     26425 => "00000010",
                     26426 => "10111001",
                     26427 => "00001110",
                     26428 => "00000010",
                     26429 => "00001001",
                     26430 => "01000000",
                     26431 => "10011001",
                     26432 => "00001110",
                     26433 => "00000010",
                     26434 => "01001100",
                     26435 => "01101011",
                     26436 => "11101011",
                     26437 => "11111100",
                     26438 => "11111100",
                     26439 => "10101010",
                     26440 => "10101011",
                     26441 => "10101100",
                     26442 => "10101101",
                     26443 => "11111100",
                     26444 => "11111100",
                     26445 => "10101110",
                     26446 => "10101111",
                     26447 => "10110000",
                     26448 => "10110001",
                     26449 => "11111100",
                     26450 => "10100101",
                     26451 => "10100110",
                     26452 => "10100111",
                     26453 => "10101000",
                     26454 => "10101001",
                     26455 => "11111100",
                     26456 => "10100000",
                     26457 => "10100001",
                     26458 => "10100010",
                     26459 => "10100011",
                     26460 => "10100100",
                     26461 => "01101001",
                     26462 => "10100101",
                     26463 => "01101010",
                     26464 => "10100111",
                     26465 => "10101000",
                     26466 => "10101001",
                     26467 => "01101011",
                     26468 => "10100000",
                     26469 => "01101100",
                     26470 => "10100010",
                     26471 => "10100011",
                     26472 => "10100100",
                     26473 => "11111100",
                     26474 => "11111100",
                     26475 => "10010110",
                     26476 => "10010111",
                     26477 => "10011000",
                     26478 => "10011001",
                     26479 => "11111100",
                     26480 => "11111100",
                     26481 => "10011010",
                     26482 => "10011011",
                     26483 => "10011100",
                     26484 => "10011101",
                     26485 => "11111100",
                     26486 => "11111100",
                     26487 => "10001111",
                     26488 => "10001110",
                     26489 => "10001110",
                     26490 => "10001111",
                     26491 => "11111100",
                     26492 => "11111100",
                     26493 => "10010101",
                     26494 => "10010100",
                     26495 => "10010100",
                     26496 => "10010101",
                     26497 => "11111100",
                     26498 => "11111100",
                     26499 => "11011100",
                     26500 => "11011100",
                     26501 => "11011111",
                     26502 => "11011111",
                     26503 => "11011100",
                     26504 => "11011100",
                     26505 => "11011101",
                     26506 => "11011101",
                     26507 => "11011110",
                     26508 => "11011110",
                     26509 => "11111100",
                     26510 => "11111100",
                     26511 => "10110010",
                     26512 => "10110011",
                     26513 => "10110100",
                     26514 => "10110101",
                     26515 => "11111100",
                     26516 => "11111100",
                     26517 => "10110110",
                     26518 => "10110011",
                     26519 => "10110111",
                     26520 => "10110101",
                     26521 => "11111100",
                     26522 => "11111100",
                     26523 => "01110000",
                     26524 => "01110001",
                     26525 => "01110010",
                     26526 => "01110011",
                     26527 => "11111100",
                     26528 => "11111100",
                     26529 => "01101110",
                     26530 => "01101110",
                     26531 => "01101111",
                     26532 => "01101111",
                     26533 => "11111100",
                     26534 => "11111100",
                     26535 => "01101101",
                     26536 => "01101101",
                     26537 => "01101111",
                     26538 => "01101111",
                     26539 => "11111100",
                     26540 => "11111100",
                     26541 => "01101111",
                     26542 => "01101111",
                     26543 => "01101110",
                     26544 => "01101110",
                     26545 => "11111100",
                     26546 => "11111100",
                     26547 => "01101111",
                     26548 => "01101111",
                     26549 => "01101101",
                     26550 => "01101101",
                     26551 => "11111100",
                     26552 => "11111100",
                     26553 => "11110100",
                     26554 => "11110100",
                     26555 => "11110101",
                     26556 => "11110101",
                     26557 => "11111100",
                     26558 => "11111100",
                     26559 => "11110100",
                     26560 => "11110100",
                     26561 => "11110101",
                     26562 => "11110101",
                     26563 => "11111100",
                     26564 => "11111100",
                     26565 => "11110101",
                     26566 => "11110101",
                     26567 => "11110100",
                     26568 => "11110100",
                     26569 => "11111100",
                     26570 => "11111100",
                     26571 => "11110101",
                     26572 => "11110101",
                     26573 => "11110100",
                     26574 => "11110100",
                     26575 => "11111100",
                     26576 => "11111100",
                     26577 => "11111100",
                     26578 => "11111100",
                     26579 => "11101111",
                     26580 => "11101111",
                     26581 => "10111001",
                     26582 => "10111000",
                     26583 => "10111011",
                     26584 => "10111010",
                     26585 => "10111100",
                     26586 => "10111100",
                     26587 => "11111100",
                     26588 => "11111100",
                     26589 => "10111101",
                     26590 => "10111101",
                     26591 => "10111100",
                     26592 => "10111100",
                     26593 => "01111010",
                     26594 => "01111011",
                     26595 => "11011010",
                     26596 => "11011011",
                     26597 => "11011000",
                     26598 => "11011000",
                     26599 => "11001101",
                     26600 => "11001101",
                     26601 => "11001110",
                     26602 => "11001110",
                     26603 => "11001111",
                     26604 => "11001111",
                     26605 => "01111101",
                     26606 => "01111100",
                     26607 => "11010001",
                     26608 => "10001100",
                     26609 => "11010011",
                     26610 => "11010010",
                     26611 => "01111101",
                     26612 => "01111100",
                     26613 => "10001001",
                     26614 => "10001000",
                     26615 => "10001011",
                     26616 => "10001010",
                     26617 => "11010101",
                     26618 => "11010100",
                     26619 => "11100011",
                     26620 => "11100010",
                     26621 => "11010011",
                     26622 => "11010010",
                     26623 => "11010101",
                     26624 => "11010100",
                     26625 => "11100011",
                     26626 => "11100010",
                     26627 => "10001011",
                     26628 => "10001010",
                     26629 => "11100101",
                     26630 => "11100101",
                     26631 => "11100110",
                     26632 => "11100110",
                     26633 => "11101011",
                     26634 => "11101011",
                     26635 => "11101100",
                     26636 => "11101100",
                     26637 => "11101101",
                     26638 => "11101101",
                     26639 => "11101110",
                     26640 => "11101110",
                     26641 => "11111100",
                     26642 => "11111100",
                     26643 => "11010000",
                     26644 => "11010000",
                     26645 => "11010111",
                     26646 => "11010111",
                     26647 => "10111111",
                     26648 => "10111110",
                     26649 => "11000001",
                     26650 => "11000000",
                     26651 => "11000010",
                     26652 => "11111100",
                     26653 => "11000100",
                     26654 => "11000011",
                     26655 => "11000110",
                     26656 => "11000101",
                     26657 => "11001000",
                     26658 => "11000111",
                     26659 => "10111111",
                     26660 => "10111110",
                     26661 => "11001010",
                     26662 => "11001001",
                     26663 => "11000010",
                     26664 => "11111100",
                     26665 => "11000100",
                     26666 => "11000011",
                     26667 => "11000110",
                     26668 => "11000101",
                     26669 => "11001100",
                     26670 => "11001011",
                     26671 => "11111100",
                     26672 => "11111100",
                     26673 => "11101000",
                     26674 => "11100111",
                     26675 => "11101010",
                     26676 => "11101001",
                     26677 => "11110010",
                     26678 => "11110010",
                     26679 => "11110011",
                     26680 => "11110011",
                     26681 => "11110010",
                     26682 => "11110010",
                     26683 => "11110001",
                     26684 => "11110001",
                     26685 => "11110001",
                     26686 => "11110001",
                     26687 => "11111100",
                     26688 => "11111100",
                     26689 => "11110000",
                     26690 => "11110000",
                     26691 => "11111100",
                     26692 => "11111100",
                     26693 => "11111100",
                     26694 => "11111100",
                     26695 => "00001100",
                     26696 => "00001100",
                     26697 => "00000000",
                     26698 => "00001100",
                     26699 => "00001100",
                     26700 => "10101000",
                     26701 => "01010100",
                     26702 => "00111100",
                     26703 => "11101010",
                     26704 => "00011000",
                     26705 => "01001000",
                     26706 => "01001000",
                     26707 => "11001100",
                     26708 => "11000000",
                     26709 => "00011000",
                     26710 => "00011000",
                     26711 => "00011000",
                     26712 => "10010000",
                     26713 => "00100100",
                     26714 => "11111111",
                     26715 => "01001000",
                     26716 => "10011100",
                     26717 => "11010010",
                     26718 => "11011000",
                     26719 => "11110000",
                     26720 => "11110110",
                     26721 => "11111100",
                     26722 => "00000001",
                     26723 => "00000010",
                     26724 => "00000011",
                     26725 => "00000010",
                     26726 => "00000001",
                     26727 => "00000001",
                     26728 => "00000011",
                     26729 => "00000011",
                     26730 => "00000011",
                     26731 => "00000001",
                     26732 => "00000001",
                     26733 => "00000010",
                     26734 => "00000010",
                     26735 => "00100001",
                     26736 => "00000001",
                     26737 => "00000010",
                     26738 => "00000001",
                     26739 => "00000001",
                     26740 => "00000010",
                     26741 => "11111111",
                     26742 => "00000010",
                     26743 => "00000010",
                     26744 => "00000001",
                     26745 => "00000001",
                     26746 => "00000010",
                     26747 => "00000010",
                     26748 => "00000010",
                     26749 => "00001000",
                     26750 => "00011000",
                     26751 => "00011000",
                     26752 => "00011001",
                     26753 => "00011010",
                     26754 => "00011001",
                     26755 => "00011000",
                     26756 => "10110101",
                     26757 => "11001111",
                     26758 => "10000101",
                     26759 => "00000010",
                     26760 => "10101101",
                     26761 => "10101110",
                     26762 => "00000011",
                     26763 => "10000101",
                     26764 => "00000101",
                     26765 => "10111100",
                     26766 => "11100101",
                     26767 => "00000110",
                     26768 => "10000100",
                     26769 => "11101011",
                     26770 => "10101001",
                     26771 => "00000000",
                     26772 => "10001101",
                     26773 => "00001001",
                     26774 => "00000001",
                     26775 => "10110101",
                     26776 => "01000110",
                     26777 => "10000101",
                     26778 => "00000011",
                     26779 => "10111101",
                     26780 => "11000101",
                     26781 => "00000011",
                     26782 => "10000101",
                     26783 => "00000100",
                     26784 => "10110101",
                     26785 => "00010110",
                     26786 => "11001001",
                     26787 => "00001101",
                     26788 => "11010000",
                     26789 => "00001010",
                     26790 => "10110100",
                     26791 => "01011000",
                     26792 => "00110000",
                     26793 => "00000110",
                     26794 => "10111100",
                     26795 => "10001010",
                     26796 => "00000111",
                     26797 => "11110000",
                     26798 => "00000001",
                     26799 => "01100000",
                     26800 => "10110101",
                     26801 => "00011110",
                     26802 => "10000101",
                     26803 => "11101101",
                     26804 => "00101001",
                     26805 => "00011111",
                     26806 => "10101000",
                     26807 => "10110101",
                     26808 => "00010110",
                     26809 => "11001001",
                     26810 => "00110101",
                     26811 => "11010000",
                     26812 => "00001000",
                     26813 => "10100000",
                     26814 => "00000000",
                     26815 => "10101001",
                     26816 => "00000001",
                     26817 => "10000101",
                     26818 => "00000011",
                     26819 => "10101001",
                     26820 => "00010101",
                     26821 => "11001001",
                     26822 => "00110011",
                     26823 => "11010000",
                     26824 => "00010011",
                     26825 => "11000110",
                     26826 => "00000010",
                     26827 => "10101001",
                     26828 => "00000011",
                     26829 => "10111100",
                     26830 => "10001010",
                     26831 => "00000111",
                     26832 => "11110000",
                     26833 => "00000010",
                     26834 => "00001001",
                     26835 => "00100000",
                     26836 => "10000101",
                     26837 => "00000100",
                     26838 => "10100000",
                     26839 => "00000000",
                     26840 => "10000100",
                     26841 => "11101101",
                     26842 => "10101001",
                     26843 => "00001000",
                     26844 => "11001001",
                     26845 => "00110010",
                     26846 => "11010000",
                     26847 => "00001000",
                     26848 => "10100000",
                     26849 => "00000011",
                     26850 => "10101110",
                     26851 => "00001110",
                     26852 => "00000111",
                     26853 => "10111101",
                     26854 => "01111111",
                     26855 => "11101000",
                     26856 => "10000101",
                     26857 => "11101111",
                     26858 => "10000100",
                     26859 => "11101100",
                     26860 => "10100110",
                     26861 => "00001000",
                     26862 => "11001001",
                     26863 => "00001100",
                     26864 => "11010000",
                     26865 => "00000111",
                     26866 => "10110101",
                     26867 => "10100000",
                     26868 => "00110000",
                     26869 => "00000011",
                     26870 => "11101110",
                     26871 => "00001001",
                     26872 => "00000001",
                     26873 => "10101101",
                     26874 => "01101010",
                     26875 => "00000011",
                     26876 => "11110000",
                     26877 => "00001001",
                     26878 => "10100000",
                     26879 => "00010110",
                     26880 => "11001001",
                     26881 => "00000001",
                     26882 => "11110000",
                     26883 => "00000001",
                     26884 => "11001000",
                     26885 => "10000100",
                     26886 => "11101111",
                     26887 => "10100100",
                     26888 => "11101111",
                     26889 => "11000000",
                     26890 => "00000110",
                     26891 => "11010000",
                     26892 => "00011101",
                     26893 => "10110101",
                     26894 => "00011110",
                     26895 => "11001001",
                     26896 => "00000010",
                     26897 => "10010000",
                     26898 => "00000100",
                     26899 => "10100010",
                     26900 => "00000100",
                     26901 => "10000110",
                     26902 => "11101100",
                     26903 => "00101001",
                     26904 => "00100000",
                     26905 => "00001101",
                     26906 => "01000111",
                     26907 => "00000111",
                     26908 => "11010000",
                     26909 => "00001100",
                     26910 => "10100101",
                     26911 => "00001001",
                     26912 => "00101001",
                     26913 => "00001000",
                     26914 => "11010000",
                     26915 => "00000110",
                     26916 => "10100101",
                     26917 => "00000011",
                     26918 => "01001001",
                     26919 => "00000011",
                     26920 => "10000101",
                     26921 => "00000011",
                     26922 => "10111001",
                     26923 => "01100010",
                     26924 => "11101000",
                     26925 => "00000101",
                     26926 => "00000100",
                     26927 => "10000101",
                     26928 => "00000100",
                     26929 => "10111001",
                     26930 => "01000111",
                     26931 => "11101000",
                     26932 => "10101010",
                     26933 => "10100100",
                     26934 => "11101100",
                     26935 => "10101101",
                     26936 => "01101010",
                     26937 => "00000011",
                     26938 => "11110000",
                     26939 => "00110000",
                     26940 => "11001001",
                     26941 => "00000001",
                     26942 => "11010000",
                     26943 => "00010011",
                     26944 => "10101101",
                     26945 => "01100011",
                     26946 => "00000011",
                     26947 => "00010000",
                     26948 => "00000010",
                     26949 => "10100010",
                     26950 => "11011110",
                     26951 => "10100101",
                     26952 => "11101101",
                     26953 => "00101001",
                     26954 => "00100000",
                     26955 => "11110000",
                     26956 => "00000011",
                     26957 => "10001110",
                     26958 => "00001001",
                     26959 => "00000001",
                     26960 => "01001100",
                     26961 => "01010010",
                     26962 => "11101010",
                     26963 => "10101101",
                     26964 => "01100011",
                     26965 => "00000011",
                     26966 => "00101001",
                     26967 => "00000001",
                     26968 => "11110000",
                     26969 => "00000010",
                     26970 => "10100010",
                     26971 => "11100100",
                     26972 => "10100101",
                     26973 => "11101101",
                     26974 => "00101001",
                     26975 => "00100000",
                     26976 => "11110000",
                     26977 => "11101110",
                     26978 => "10100101",
                     26979 => "00000010",
                     26980 => "00111000",
                     26981 => "11101001",
                     26982 => "00010000",
                     26983 => "10000101",
                     26984 => "00000010",
                     26985 => "01001100",
                     26986 => "01001101",
                     26987 => "11101001",
                     26988 => "11100000",
                     26989 => "00100100",
                     26990 => "11010000",
                     26991 => "00010001",
                     26992 => "11000000",
                     26993 => "00000101",
                     26994 => "11010000",
                     26995 => "00001010",
                     26996 => "10100010",
                     26997 => "00110000",
                     26998 => "10101001",
                     26999 => "00000010",
                     27000 => "10000101",
                     27001 => "00000011",
                     27002 => "10101001",
                     27003 => "00000101",
                     27004 => "10000101",
                     27005 => "11101100",
                     27006 => "01001100",
                     27007 => "11010001",
                     27008 => "11101001",
                     27009 => "11100000",
                     27010 => "10010000",
                     27011 => "11010000",
                     27012 => "00010010",
                     27013 => "10100101",
                     27014 => "11101101",
                     27015 => "00101001",
                     27016 => "00100000",
                     27017 => "11010000",
                     27018 => "00001001",
                     27019 => "10101101",
                     27020 => "10001111",
                     27021 => "00000111",
                     27022 => "11001001",
                     27023 => "00010000",
                     27024 => "10110000",
                     27025 => "00000010",
                     27026 => "10100010",
                     27027 => "10010110",
                     27028 => "01001100",
                     27029 => "00111110",
                     27030 => "11101010",
                     27031 => "10100101",
                     27032 => "11101111",
                     27033 => "11001001",
                     27034 => "00000100",
                     27035 => "10110000",
                     27036 => "00010000",
                     27037 => "11000000",
                     27038 => "00000010",
                     27039 => "10010000",
                     27040 => "00001100",
                     27041 => "10100010",
                     27042 => "01011010",
                     27043 => "10100100",
                     27044 => "11101111",
                     27045 => "11000000",
                     27046 => "00000010",
                     27047 => "11010000",
                     27048 => "00000100",
                     27049 => "10100010",
                     27050 => "01111110",
                     27051 => "11100110",
                     27052 => "00000010",
                     27053 => "10100101",
                     27054 => "11101100",
                     27055 => "11001001",
                     27056 => "00000100",
                     27057 => "11010000",
                     27058 => "00011110",
                     27059 => "10100010",
                     27060 => "01110010",
                     27061 => "11100110",
                     27062 => "00000010",
                     27063 => "10100100",
                     27064 => "11101111",
                     27065 => "11000000",
                     27066 => "00000010",
                     27067 => "11110000",
                     27068 => "00000100",
                     27069 => "10100010",
                     27070 => "01100110",
                     27071 => "11100110",
                     27072 => "00000010",
                     27073 => "11000000",
                     27074 => "00000110",
                     27075 => "11010000",
                     27076 => "00001100",
                     27077 => "10100010",
                     27078 => "01010100",
                     27079 => "10100101",
                     27080 => "11101101",
                     27081 => "00101001",
                     27082 => "00100000",
                     27083 => "11010000",
                     27084 => "00000100",
                     27085 => "10100010",
                     27086 => "10001010",
                     27087 => "11000110",
                     27088 => "00000010",
                     27089 => "10100100",
                     27090 => "00001000",
                     27091 => "10100101",
                     27092 => "11101111",
                     27093 => "11001001",
                     27094 => "00000101",
                     27095 => "11010000",
                     27096 => "00001100",
                     27097 => "10100101",
                     27098 => "11101101",
                     27099 => "11110000",
                     27100 => "00100100",
                     27101 => "00101001",
                     27102 => "00001000",
                     27103 => "11110000",
                     27104 => "01011101",
                     27105 => "10100010",
                     27106 => "10110100",
                     27107 => "11010000",
                     27108 => "00011100",
                     27109 => "11100000",
                     27110 => "01001000",
                     27111 => "11110000",
                     27112 => "00011000",
                     27113 => "10111001",
                     27114 => "10010110",
                     27115 => "00000111",
                     27116 => "11001001",
                     27117 => "00000101",
                     27118 => "10110000",
                     27119 => "01001110",
                     27120 => "11100000",
                     27121 => "00111100",
                     27122 => "11010000",
                     27123 => "00001101",
                     27124 => "11001001",
                     27125 => "00000001",
                     27126 => "11110000",
                     27127 => "01000110",
                     27128 => "11100110",
                     27129 => "00000010",
                     27130 => "11100110",
                     27131 => "00000010",
                     27132 => "11100110",
                     27133 => "00000010",
                     27134 => "01001100",
                     27135 => "00110000",
                     27136 => "11101010",
                     27137 => "10100101",
                     27138 => "11101111",
                     27139 => "11001001",
                     27140 => "00000110",
                     27141 => "11110000",
                     27142 => "00110111",
                     27143 => "11001001",
                     27144 => "00001000",
                     27145 => "11110000",
                     27146 => "00110011",
                     27147 => "11001001",
                     27148 => "00001100",
                     27149 => "11110000",
                     27150 => "00101111",
                     27151 => "11001001",
                     27152 => "00011000",
                     27153 => "10110000",
                     27154 => "00101011",
                     27155 => "10100000",
                     27156 => "00000000",
                     27157 => "11001001",
                     27158 => "00010101",
                     27159 => "11010000",
                     27160 => "00010000",
                     27161 => "11001000",
                     27162 => "10101101",
                     27163 => "01011111",
                     27164 => "00000111",
                     27165 => "11001001",
                     27166 => "00000111",
                     27167 => "10110000",
                     27168 => "00011101",
                     27169 => "10100010",
                     27170 => "10100010",
                     27171 => "10101001",
                     27172 => "00000011",
                     27173 => "10000101",
                     27174 => "11101100",
                     27175 => "11010000",
                     27176 => "00010101",
                     27177 => "10100101",
                     27178 => "00001001",
                     27179 => "00111001",
                     27180 => "01111101",
                     27181 => "11101000",
                     27182 => "11010000",
                     27183 => "00001110",
                     27184 => "10100101",
                     27185 => "11101101",
                     27186 => "00101001",
                     27187 => "10100000",
                     27188 => "00001101",
                     27189 => "01000111",
                     27190 => "00000111",
                     27191 => "11010000",
                     27192 => "00000101",
                     27193 => "10001010",
                     27194 => "00011000",
                     27195 => "01101001",
                     27196 => "00000110",
                     27197 => "10101010",
                     27198 => "10100101",
                     27199 => "11101101",
                     27200 => "00101001",
                     27201 => "00100000",
                     27202 => "11110000",
                     27203 => "00001110",
                     27204 => "10100101",
                     27205 => "11101111",
                     27206 => "11001001",
                     27207 => "00000100",
                     27208 => "10010000",
                     27209 => "00001000",
                     27210 => "10100000",
                     27211 => "00000001",
                     27212 => "10001100",
                     27213 => "00001001",
                     27214 => "00000001",
                     27215 => "10001000",
                     27216 => "10000100",
                     27217 => "11101100",
                     27218 => "10100100",
                     27219 => "11101011",
                     27220 => "00100000",
                     27221 => "10110001",
                     27222 => "11101011",
                     27223 => "00100000",
                     27224 => "10110001",
                     27225 => "11101011",
                     27226 => "00100000",
                     27227 => "10110001",
                     27228 => "11101011",
                     27229 => "10100110",
                     27230 => "00001000",
                     27231 => "10111100",
                     27232 => "11100101",
                     27233 => "00000110",
                     27234 => "10100101",
                     27235 => "11101111",
                     27236 => "11001001",
                     27237 => "00001000",
                     27238 => "11010000",
                     27239 => "00000011",
                     27240 => "01001100",
                     27241 => "01101011",
                     27242 => "11101011",
                     27243 => "10101101",
                     27244 => "00001001",
                     27245 => "00000001",
                     27246 => "11110000",
                     27247 => "00111101",
                     27248 => "10111001",
                     27249 => "00000010",
                     27250 => "00000010",
                     27251 => "00001001",
                     27252 => "10000000",
                     27253 => "11001000",
                     27254 => "11001000",
                     27255 => "00100000",
                     27256 => "10111100",
                     27257 => "11100101",
                     27258 => "10001000",
                     27259 => "10001000",
                     27260 => "10011000",
                     27261 => "10101010",
                     27262 => "10100101",
                     27263 => "11101111",
                     27264 => "11001001",
                     27265 => "00000101",
                     27266 => "11110000",
                     27267 => "00001101",
                     27268 => "11001001",
                     27269 => "00010001",
                     27270 => "11110000",
                     27271 => "00001001",
                     27272 => "11001001",
                     27273 => "00010101",
                     27274 => "10110000",
                     27275 => "00000101",
                     27276 => "10001010",
                     27277 => "00011000",
                     27278 => "01101001",
                     27279 => "00001000",
                     27280 => "10101010",
                     27281 => "10111101",
                     27282 => "00000001",
                     27283 => "00000010",
                     27284 => "01001000",
                     27285 => "10111101",
                     27286 => "00000101",
                     27287 => "00000010",
                     27288 => "01001000",
                     27289 => "10111001",
                     27290 => "00010001",
                     27291 => "00000010",
                     27292 => "10011101",
                     27293 => "00000001",
                     27294 => "00000010",
                     27295 => "10111001",
                     27296 => "00010101",
                     27297 => "00000010",
                     27298 => "10011101",
                     27299 => "00000101",
                     27300 => "00000010",
                     27301 => "01101000",
                     27302 => "10011001",
                     27303 => "00010101",
                     27304 => "00000010",
                     27305 => "01101000",
                     27306 => "10011001",
                     27307 => "00010001",
                     27308 => "00000010",
                     27309 => "10101101",
                     27310 => "01101010",
                     27311 => "00000011",
                     27312 => "11010000",
                     27313 => "10110110",
                     27314 => "10100101",
                     27315 => "11101111",
                     27316 => "10100110",
                     27317 => "11101100",
                     27318 => "11001001",
                     27319 => "00000101",
                     27320 => "11010000",
                     27321 => "00000011",
                     27322 => "01001100",
                     27323 => "01101011",
                     27324 => "11101011",
                     27325 => "11001001",
                     27326 => "00000111",
                     27327 => "11110000",
                     27328 => "00011101",
                     27329 => "11001001",
                     27330 => "00001101",
                     27331 => "11110000",
                     27332 => "00011001",
                     27333 => "11001001",
                     27334 => "00001100",
                     27335 => "11110000",
                     27336 => "00010101",
                     27337 => "11001001",
                     27338 => "00010010",
                     27339 => "11010000",
                     27340 => "00000100",
                     27341 => "11100000",
                     27342 => "00000101",
                     27343 => "11010000",
                     27344 => "01001000",
                     27345 => "11001001",
                     27346 => "00010101",
                     27347 => "11010000",
                     27348 => "00000101",
                     27349 => "10101001",
                     27350 => "01000010",
                     27351 => "10011001",
                     27352 => "00010110",
                     27353 => "00000010",
                     27354 => "11100000",
                     27355 => "00000010",
                     27356 => "10010000",
                     27357 => "00111011",
                     27358 => "10101101",
                     27359 => "01101010",
                     27360 => "00000011",
                     27361 => "11010000",
                     27362 => "00110110",
                     27363 => "10111001",
                     27364 => "00000010",
                     27365 => "00000010",
                     27366 => "00101001",
                     27367 => "10100011",
                     27368 => "10011001",
                     27369 => "00000010",
                     27370 => "00000010",
                     27371 => "10011001",
                     27372 => "00001010",
                     27373 => "00000010",
                     27374 => "10011001",
                     27375 => "00010010",
                     27376 => "00000010",
                     27377 => "00001001",
                     27378 => "01000000",
                     27379 => "11100000",
                     27380 => "00000101",
                     27381 => "11010000",
                     27382 => "00000010",
                     27383 => "00001001",
                     27384 => "10000000",
                     27385 => "10011001",
                     27386 => "00000110",
                     27387 => "00000010",
                     27388 => "10011001",
                     27389 => "00001110",
                     27390 => "00000010",
                     27391 => "10011001",
                     27392 => "00010110",
                     27393 => "00000010",
                     27394 => "11100000",
                     27395 => "00000100",
                     27396 => "11010000",
                     27397 => "00010011",
                     27398 => "10111001",
                     27399 => "00001010",
                     27400 => "00000010",
                     27401 => "00001001",
                     27402 => "10000000",
                     27403 => "10011001",
                     27404 => "00001010",
                     27405 => "00000010",
                     27406 => "10011001",
                     27407 => "00010010",
                     27408 => "00000010",
                     27409 => "00001001",
                     27410 => "01000000",
                     27411 => "10011001",
                     27412 => "00001110",
                     27413 => "00000010",
                     27414 => "10011001",
                     27415 => "00010110",
                     27416 => "00000010",
                     27417 => "10100101",
                     27418 => "11101111",
                     27419 => "11001001",
                     27420 => "00010001",
                     27421 => "11010000",
                     27422 => "00110110",
                     27423 => "10101101",
                     27424 => "00001001",
                     27425 => "00000001",
                     27426 => "11010000",
                     27427 => "00100001",
                     27428 => "10111001",
                     27429 => "00010010",
                     27430 => "00000010",
                     27431 => "00101001",
                     27432 => "10000001",
                     27433 => "10011001",
                     27434 => "00010010",
                     27435 => "00000010",
                     27436 => "10111001",
                     27437 => "00010110",
                     27438 => "00000010",
                     27439 => "00001001",
                     27440 => "01000001",
                     27441 => "10011001",
                     27442 => "00010110",
                     27443 => "00000010",
                     27444 => "10101110",
                     27445 => "10001111",
                     27446 => "00000111",
                     27447 => "11100000",
                     27448 => "00010000",
                     27449 => "10110000",
                     27450 => "00110000",
                     27451 => "10011001",
                     27452 => "00001110",
                     27453 => "00000010",
                     27454 => "00101001",
                     27455 => "10000001",
                     27456 => "10011001",
                     27457 => "00001010",
                     27458 => "00000010",
                     27459 => "10010000",
                     27460 => "00100110",
                     27461 => "10111001",
                     27462 => "00000010",
                     27463 => "00000010",
                     27464 => "00101001",
                     27465 => "10000001",
                     27466 => "10011001",
                     27467 => "00000010",
                     27468 => "00000010",
                     27469 => "10111001",
                     27470 => "00000110",
                     27471 => "00000010",
                     27472 => "00001001",
                     27473 => "01000001",
                     27474 => "10011001",
                     27475 => "00000110",
                     27476 => "00000010",
                     27477 => "10100101",
                     27478 => "11101111",
                     27479 => "11001001",
                     27480 => "00011000",
                     27481 => "10010000",
                     27482 => "00010000",
                     27483 => "10101001",
                     27484 => "10000010",
                     27485 => "10011001",
                     27486 => "00001010",
                     27487 => "00000010",
                     27488 => "10011001",
                     27489 => "00010010",
                     27490 => "00000010",
                     27491 => "00001001",
                     27492 => "01000000",
                     27493 => "10011001",
                     27494 => "00001110",
                     27495 => "00000010",
                     27496 => "10011001",
                     27497 => "00010110",
                     27498 => "00000010",
                     27499 => "10100110",
                     27500 => "00001000",
                     27501 => "10101101",
                     27502 => "11010001",
                     27503 => "00000011",
                     27504 => "01001010",
                     27505 => "01001010",
                     27506 => "01001010",
                     27507 => "01001000",
                     27508 => "10010000",
                     27509 => "00000101",
                     27510 => "10101001",
                     27511 => "00000100",
                     27512 => "00100000",
                     27513 => "11001000",
                     27514 => "11101011",
                     27515 => "01101000",
                     27516 => "01001010",
                     27517 => "01001000",
                     27518 => "10010000",
                     27519 => "00000101",
                     27520 => "10101001",
                     27521 => "00000000",
                     27522 => "00100000",
                     27523 => "11001000",
                     27524 => "11101011",
                     27525 => "01101000",
                     27526 => "01001010",
                     27527 => "01001010",
                     27528 => "01001000",
                     27529 => "10010000",
                     27530 => "00000101",
                     27531 => "10101001",
                     27532 => "00010000",
                     27533 => "00100000",
                     27534 => "10111110",
                     27535 => "11101011",
                     27536 => "01101000",
                     27537 => "01001010",
                     27538 => "01001000",
                     27539 => "10010000",
                     27540 => "00000101",
                     27541 => "10101001",
                     27542 => "00001000",
                     27543 => "00100000",
                     27544 => "10111110",
                     27545 => "11101011",
                     27546 => "01101000",
                     27547 => "01001010",
                     27548 => "10010000",
                     27549 => "00010010",
                     27550 => "00100000",
                     27551 => "10111110",
                     27552 => "11101011",
                     27553 => "10110101",
                     27554 => "00010110",
                     27555 => "11001001",
                     27556 => "00001100",
                     27557 => "11110000",
                     27558 => "00001001",
                     27559 => "10110101",
                     27560 => "10110110",
                     27561 => "11001001",
                     27562 => "00000010",
                     27563 => "11010000",
                     27564 => "00000011",
                     27565 => "00100000",
                     27566 => "10011110",
                     27567 => "11001001",
                     27568 => "01100000",
                     27569 => "10111101",
                     27570 => "01000101",
                     27571 => "11100111",
                     27572 => "10000101",
                     27573 => "00000000",
                     27574 => "10111101",
                     27575 => "01000110",
                     27576 => "11100111",
                     27577 => "10000101",
                     27578 => "00000001",
                     27579 => "01001100",
                     27580 => "10001001",
                     27581 => "11110010",
                     27582 => "00011000",
                     27583 => "01111101",
                     27584 => "11100101",
                     27585 => "00000110",
                     27586 => "10101000",
                     27587 => "10101001",
                     27588 => "11111000",
                     27589 => "01001100",
                     27590 => "11001000",
                     27591 => "11100101",
                     27592 => "00011000",
                     27593 => "01111101",
                     27594 => "11100101",
                     27595 => "00000110",
                     27596 => "10101000",
                     27597 => "00100000",
                     27598 => "01010001",
                     27599 => "11101100",
                     27600 => "10011001",
                     27601 => "00010000",
                     27602 => "00000010",
                     27603 => "01100000",
                     27604 => "10000101",
                     27605 => "10000101",
                     27606 => "10000110",
                     27607 => "10000110",
                     27608 => "10101101",
                     27609 => "10111100",
                     27610 => "00000011",
                     27611 => "10000101",
                     27612 => "00000010",
                     27613 => "10101101",
                     27614 => "10110001",
                     27615 => "00000011",
                     27616 => "10000101",
                     27617 => "00000101",
                     27618 => "10101001",
                     27619 => "00000011",
                     27620 => "10000101",
                     27621 => "00000100",
                     27622 => "01001010",
                     27623 => "10000101",
                     27624 => "00000011",
                     27625 => "10111100",
                     27626 => "11101100",
                     27627 => "00000110",
                     27628 => "10100010",
                     27629 => "00000000",
                     27630 => "10111101",
                     27631 => "11010100",
                     27632 => "11101011",
                     27633 => "10000101",
                     27634 => "00000000",
                     27635 => "10111101",
                     27636 => "11010101",
                     27637 => "11101011",
                     27638 => "00100000",
                     27639 => "10111001",
                     27640 => "11101011",
                     27641 => "11100000",
                     27642 => "00000100",
                     27643 => "11010000",
                     27644 => "11110001",
                     27645 => "10100110",
                     27646 => "00001000",
                     27647 => "10111100",
                     27648 => "11101100",
                     27649 => "00000110",
                     27650 => "10101101",
                     27651 => "01001110",
                     27652 => "00000111",
                     27653 => "11001001",
                     27654 => "00000001",
                     27655 => "11110000",
                     27656 => "00001000",
                     27657 => "10101001",
                     27658 => "10000110",
                     27659 => "10011001",
                     27660 => "00000001",
                     27661 => "00000010",
                     27662 => "10011001",
                     27663 => "00000101",
                     27664 => "00000010",
                     27665 => "10111101",
                     27666 => "11101000",
                     27667 => "00000011",
                     27668 => "11001001",
                     27669 => "11000100",
                     27670 => "11010000",
                     27671 => "00100100",
                     27672 => "10101001",
                     27673 => "10000111",
                     27674 => "11001000",
                     27675 => "00100000",
                     27676 => "11000010",
                     27677 => "11100101",
                     27678 => "10001000",
                     27679 => "10101001",
                     27680 => "00000011",
                     27681 => "10101110",
                     27682 => "01001110",
                     27683 => "00000111",
                     27684 => "11001010",
                     27685 => "11110000",
                     27686 => "00000001",
                     27687 => "01001010",
                     27688 => "10100110",
                     27689 => "00001000",
                     27690 => "10011001",
                     27691 => "00000010",
                     27692 => "00000010",
                     27693 => "00001001",
                     27694 => "01000000",
                     27695 => "10011001",
                     27696 => "00000110",
                     27697 => "00000010",
                     27698 => "00001001",
                     27699 => "10000000",
                     27700 => "10011001",
                     27701 => "00001110",
                     27702 => "00000010",
                     27703 => "00101001",
                     27704 => "10000011",
                     27705 => "10011001",
                     27706 => "00001010",
                     27707 => "00000010",
                     27708 => "10101101",
                     27709 => "11010100",
                     27710 => "00000011",
                     27711 => "01001000",
                     27712 => "00101001",
                     27713 => "00000100",
                     27714 => "11110000",
                     27715 => "00001000",
                     27716 => "10101001",
                     27717 => "11111000",
                     27718 => "10011001",
                     27719 => "00000100",
                     27720 => "00000010",
                     27721 => "10011001",
                     27722 => "00001100",
                     27723 => "00000010",
                     27724 => "01101000",
                     27725 => "00101001",
                     27726 => "00001000",
                     27727 => "11110000",
                     27728 => "00001000",
                     27729 => "10101001",
                     27730 => "11111000",
                     27731 => "10011001",
                     27732 => "00000000",
                     27733 => "00000010",
                     27734 => "10011001",
                     27735 => "00001000",
                     27736 => "00000010",
                     27737 => "01100000",
                     27738 => "10101001",
                     27739 => "00000010",
                     27740 => "10000101",
                     27741 => "00000000",
                     27742 => "10101001",
                     27743 => "01110101",
                     27744 => "10100100",
                     27745 => "00001110",
                     27746 => "11000000",
                     27747 => "00000101",
                     27748 => "11110000",
                     27749 => "00000110",
                     27750 => "10101001",
                     27751 => "00000011",
                     27752 => "10000101",
                     27753 => "00000000",
                     27754 => "10101001",
                     27755 => "10000100",
                     27756 => "10111100",
                     27757 => "11101100",
                     27758 => "00000110",
                     27759 => "11001000",
                     27760 => "00100000",
                     27761 => "11000010",
                     27762 => "11100101",
                     27763 => "10100101",
                     27764 => "00001001",
                     27765 => "00001010",
                     27766 => "00001010",
                     27767 => "00001010",
                     27768 => "00001010",
                     27769 => "00101001",
                     27770 => "11000000",
                     27771 => "00000101",
                     27772 => "00000000",
                     27773 => "11001000",
                     27774 => "00100000",
                     27775 => "11000010",
                     27776 => "11100101",
                     27777 => "10001000",
                     27778 => "10001000",
                     27779 => "10101101",
                     27780 => "10111100",
                     27781 => "00000011",
                     27782 => "00100000",
                     27783 => "11001000",
                     27784 => "11100101",
                     27785 => "10101101",
                     27786 => "10110001",
                     27787 => "00000011",
                     27788 => "10011001",
                     27789 => "00000011",
                     27790 => "00000010",
                     27791 => "10111101",
                     27792 => "11110001",
                     27793 => "00000011",
                     27794 => "00111000",
                     27795 => "11101101",
                     27796 => "00011100",
                     27797 => "00000111",
                     27798 => "10000101",
                     27799 => "00000000",
                     27800 => "00111000",
                     27801 => "11101101",
                     27802 => "10110001",
                     27803 => "00000011",
                     27804 => "01100101",
                     27805 => "00000000",
                     27806 => "01101001",
                     27807 => "00000110",
                     27808 => "10011001",
                     27809 => "00000111",
                     27810 => "00000010",
                     27811 => "10101101",
                     27812 => "10111101",
                     27813 => "00000011",
                     27814 => "10011001",
                     27815 => "00001000",
                     27816 => "00000010",
                     27817 => "10011001",
                     27818 => "00001100",
                     27819 => "00000010",
                     27820 => "10101101",
                     27821 => "10110010",
                     27822 => "00000011",
                     27823 => "10011001",
                     27824 => "00001011",
                     27825 => "00000010",
                     27826 => "10100101",
                     27827 => "00000000",
                     27828 => "00111000",
                     27829 => "11101101",
                     27830 => "10110010",
                     27831 => "00000011",
                     27832 => "01100101",
                     27833 => "00000000",
                     27834 => "01101001",
                     27835 => "00000110",
                     27836 => "10011001",
                     27837 => "00001111",
                     27838 => "00000010",
                     27839 => "10101101",
                     27840 => "11010100",
                     27841 => "00000011",
                     27842 => "00100000",
                     27843 => "01001101",
                     27844 => "11101100",
                     27845 => "10101101",
                     27846 => "11010100",
                     27847 => "00000011",
                     27848 => "00001010",
                     27849 => "10010000",
                     27850 => "00000101",
                     27851 => "10101001",
                     27852 => "11111000",
                     27853 => "00100000",
                     27854 => "11001000",
                     27855 => "11100101",
                     27856 => "10100101",
                     27857 => "00000000",
                     27858 => "00010000",
                     27859 => "00010000",
                     27860 => "10111001",
                     27861 => "00000011",
                     27862 => "00000010",
                     27863 => "11011001",
                     27864 => "00000111",
                     27865 => "00000010",
                     27866 => "10010000",
                     27867 => "00001000",
                     27868 => "10101001",
                     27869 => "11111000",
                     27870 => "10011001",
                     27871 => "00000100",
                     27872 => "00000010",
                     27873 => "10011001",
                     27874 => "00001100",
                     27875 => "00000010",
                     27876 => "01100000",
                     27877 => "10111100",
                     27878 => "11110001",
                     27879 => "00000110",
                     27880 => "10101101",
                     27881 => "10111010",
                     27882 => "00000011",
                     27883 => "10011001",
                     27884 => "00000000",
                     27885 => "00000010",
                     27886 => "10101101",
                     27887 => "10101111",
                     27888 => "00000011",
                     27889 => "10011001",
                     27890 => "00000011",
                     27891 => "00000010",
                     27892 => "10100101",
                     27893 => "00001001",
                     27894 => "01001010",
                     27895 => "01001010",
                     27896 => "01001000",
                     27897 => "00101001",
                     27898 => "00000001",
                     27899 => "01001001",
                     27900 => "01100100",
                     27901 => "10011001",
                     27902 => "00000001",
                     27903 => "00000010",
                     27904 => "01101000",
                     27905 => "01001010",
                     27906 => "01001010",
                     27907 => "10101001",
                     27908 => "00000010",
                     27909 => "10010000",
                     27910 => "00000010",
                     27911 => "00001001",
                     27912 => "11000000",
                     27913 => "10011001",
                     27914 => "00000010",
                     27915 => "00000010",
                     27916 => "01100000",
                     27917 => "01101000",
                     27918 => "01100111",
                     27919 => "01100110",
                     27920 => "10111100",
                     27921 => "11101100",
                     27922 => "00000110",
                     27923 => "10110101",
                     27924 => "00100100",
                     27925 => "11110110",
                     27926 => "00100100",
                     27927 => "01001010",
                     27928 => "00101001",
                     27929 => "00000111",
                     27930 => "11001001",
                     27931 => "00000011",
                     27932 => "10110000",
                     27933 => "01001010",
                     27934 => "10101010",
                     27935 => "10111101",
                     27936 => "00001101",
                     27937 => "11101101",
                     27938 => "11001000",
                     27939 => "00100000",
                     27940 => "11000010",
                     27941 => "11100101",
                     27942 => "10001000",
                     27943 => "10100110",
                     27944 => "00001000",
                     27945 => "10101101",
                     27946 => "10111010",
                     27947 => "00000011",
                     27948 => "00111000",
                     27949 => "11101001",
                     27950 => "00000100",
                     27951 => "10011001",
                     27952 => "00000000",
                     27953 => "00000010",
                     27954 => "10011001",
                     27955 => "00001000",
                     27956 => "00000010",
                     27957 => "00011000",
                     27958 => "01101001",
                     27959 => "00001000",
                     27960 => "10011001",
                     27961 => "00000100",
                     27962 => "00000010",
                     27963 => "10011001",
                     27964 => "00001100",
                     27965 => "00000010",
                     27966 => "10101101",
                     27967 => "10101111",
                     27968 => "00000011",
                     27969 => "00111000",
                     27970 => "11101001",
                     27971 => "00000100",
                     27972 => "10011001",
                     27973 => "00000011",
                     27974 => "00000010",
                     27975 => "10011001",
                     27976 => "00000111",
                     27977 => "00000010",
                     27978 => "00011000",
                     27979 => "01101001",
                     27980 => "00001000",
                     27981 => "10011001",
                     27982 => "00001011",
                     27983 => "00000010",
                     27984 => "10011001",
                     27985 => "00001111",
                     27986 => "00000010",
                     27987 => "10101001",
                     27988 => "00000010",
                     27989 => "10011001",
                     27990 => "00000010",
                     27991 => "00000010",
                     27992 => "10101001",
                     27993 => "10000010",
                     27994 => "10011001",
                     27995 => "00000110",
                     27996 => "00000010",
                     27997 => "10101001",
                     27998 => "01000010",
                     27999 => "10011001",
                     28000 => "00001010",
                     28001 => "00000010",
                     28002 => "10101001",
                     28003 => "11000010",
                     28004 => "10011001",
                     28005 => "00001110",
                     28006 => "00000010",
                     28007 => "01100000",
                     28008 => "10101001",
                     28009 => "00000000",
                     28010 => "10010101",
                     28011 => "00100100",
                     28012 => "01100000",
                     28013 => "10111100",
                     28014 => "11100101",
                     28015 => "00000110",
                     28016 => "10101001",
                     28017 => "01011011",
                     28018 => "11001000",
                     28019 => "00100000",
                     28020 => "10111100",
                     28021 => "11100101",
                     28022 => "11001000",
                     28023 => "10101001",
                     28024 => "00000010",
                     28025 => "00100000",
                     28026 => "10111100",
                     28027 => "11100101",
                     28028 => "10001000",
                     28029 => "10001000",
                     28030 => "10101101",
                     28031 => "10101110",
                     28032 => "00000011",
                     28033 => "10011001",
                     28034 => "00000011",
                     28035 => "00000010",
                     28036 => "10011001",
                     28037 => "00001111",
                     28038 => "00000010",
                     28039 => "00011000",
                     28040 => "01101001",
                     28041 => "00001000",
                     28042 => "10011001",
                     28043 => "00000111",
                     28044 => "00000010",
                     28045 => "10011001",
                     28046 => "00010011",
                     28047 => "00000010",
                     28048 => "00011000",
                     28049 => "01101001",
                     28050 => "00001000",
                     28051 => "10011001",
                     28052 => "00001011",
                     28053 => "00000010",
                     28054 => "10011001",
                     28055 => "00010111",
                     28056 => "00000010",
                     28057 => "10110101",
                     28058 => "11001111",
                     28059 => "10101010",
                     28060 => "01001000",
                     28061 => "11100000",
                     28062 => "00100000",
                     28063 => "10110000",
                     28064 => "00000010",
                     28065 => "10101001",
                     28066 => "11111000",
                     28067 => "00100000",
                     28068 => "11000101",
                     28069 => "11100101",
                     28070 => "01101000",
                     28071 => "00011000",
                     28072 => "01101001",
                     28073 => "10000000",
                     28074 => "10101010",
                     28075 => "11100000",
                     28076 => "00100000",
                     28077 => "10110000",
                     28078 => "00000010",
                     28079 => "10101001",
                     28080 => "11111000",
                     28081 => "10011001",
                     28082 => "00001100",
                     28083 => "00000010",
                     28084 => "10011001",
                     28085 => "00010000",
                     28086 => "00000010",
                     28087 => "10011001",
                     28088 => "00010100",
                     28089 => "00000010",
                     28090 => "10101101",
                     28091 => "11010001",
                     28092 => "00000011",
                     28093 => "01001000",
                     28094 => "00101001",
                     28095 => "00001000",
                     28096 => "11110000",
                     28097 => "00001000",
                     28098 => "10101001",
                     28099 => "11111000",
                     28100 => "10011001",
                     28101 => "00000000",
                     28102 => "00000010",
                     28103 => "10011001",
                     28104 => "00001100",
                     28105 => "00000010",
                     28106 => "01101000",
                     28107 => "01001000",
                     28108 => "00101001",
                     28109 => "00000100",
                     28110 => "11110000",
                     28111 => "00001000",
                     28112 => "10101001",
                     28113 => "11111000",
                     28114 => "10011001",
                     28115 => "00000100",
                     28116 => "00000010",
                     28117 => "10011001",
                     28118 => "00010000",
                     28119 => "00000010",
                     28120 => "01101000",
                     28121 => "00101001",
                     28122 => "00000010",
                     28123 => "11110000",
                     28124 => "00001000",
                     28125 => "10101001",
                     28126 => "11111000",
                     28127 => "10011001",
                     28128 => "00001000",
                     28129 => "00000010",
                     28130 => "10011001",
                     28131 => "00010100",
                     28132 => "00000010",
                     28133 => "10100110",
                     28134 => "00001000",
                     28135 => "01100000",
                     28136 => "10100100",
                     28137 => "10110101",
                     28138 => "10001000",
                     28139 => "11010000",
                     28140 => "00100000",
                     28141 => "10101101",
                     28142 => "11010011",
                     28143 => "00000011",
                     28144 => "00101001",
                     28145 => "00001000",
                     28146 => "11010000",
                     28147 => "00011001",
                     28148 => "10111100",
                     28149 => "11101110",
                     28150 => "00000110",
                     28151 => "10101101",
                     28152 => "10110000",
                     28153 => "00000011",
                     28154 => "10011001",
                     28155 => "00000011",
                     28156 => "00000010",
                     28157 => "10101101",
                     28158 => "10111011",
                     28159 => "00000011",
                     28160 => "10011001",
                     28161 => "00000000",
                     28162 => "00000010",
                     28163 => "10101001",
                     28164 => "01110100",
                     28165 => "10011001",
                     28166 => "00000001",
                     28167 => "00000010",
                     28168 => "10101001",
                     28169 => "00000010",
                     28170 => "10011001",
                     28171 => "00000010",
                     28172 => "00000010",
                     28173 => "01100000",
                     28174 => "00100000",
                     28175 => "00101000",
                     28176 => "11001000",
                     28177 => "00011000",
                     28178 => "00000000",
                     28179 => "01000000",
                     28180 => "01010000",
                     28181 => "01011000",
                     28182 => "10000000",
                     28183 => "10001000",
                     28184 => "10111000",
                     28185 => "01111000",
                     28186 => "01100000",
                     28187 => "10100000",
                     28188 => "10110000",
                     28189 => "10111000",
                     28190 => "00000000",
                     28191 => "00000001",
                     28192 => "00000010",
                     28193 => "00000011",
                     28194 => "00000100",
                     28195 => "00000101",
                     28196 => "00000110",
                     28197 => "00000111",
                     28198 => "00001000",
                     28199 => "00001001",
                     28200 => "00001010",
                     28201 => "00001011",
                     28202 => "00001100",
                     28203 => "00001101",
                     28204 => "00001110",
                     28205 => "00001111",
                     28206 => "00010000",
                     28207 => "00010001",
                     28208 => "00010010",
                     28209 => "00010011",
                     28210 => "00010100",
                     28211 => "00010101",
                     28212 => "00010110",
                     28213 => "00010111",
                     28214 => "00011000",
                     28215 => "00011001",
                     28216 => "00011010",
                     28217 => "00011011",
                     28218 => "00011100",
                     28219 => "00011101",
                     28220 => "00011110",
                     28221 => "00011111",
                     28222 => "00100000",
                     28223 => "00100001",
                     28224 => "00100010",
                     28225 => "00100011",
                     28226 => "00100100",
                     28227 => "00100101",
                     28228 => "00100110",
                     28229 => "00100111",
                     28230 => "00001000",
                     28231 => "00001001",
                     28232 => "00101000",
                     28233 => "00101001",
                     28234 => "00101010",
                     28235 => "00101011",
                     28236 => "00101100",
                     28237 => "00101101",
                     28238 => "00001000",
                     28239 => "00001001",
                     28240 => "00001010",
                     28241 => "00001011",
                     28242 => "00001100",
                     28243 => "00110000",
                     28244 => "00101100",
                     28245 => "00101101",
                     28246 => "00001000",
                     28247 => "00001001",
                     28248 => "00001010",
                     28249 => "00001011",
                     28250 => "00101110",
                     28251 => "00101111",
                     28252 => "00101100",
                     28253 => "00101101",
                     28254 => "00001000",
                     28255 => "00001001",
                     28256 => "00101000",
                     28257 => "00101001",
                     28258 => "00101010",
                     28259 => "00101011",
                     28260 => "01011100",
                     28261 => "01011101",
                     28262 => "00001000",
                     28263 => "00001001",
                     28264 => "00001010",
                     28265 => "00001011",
                     28266 => "00001100",
                     28267 => "00001101",
                     28268 => "01011110",
                     28269 => "01011111",
                     28270 => "11111100",
                     28271 => "11111100",
                     28272 => "00001000",
                     28273 => "00001001",
                     28274 => "01011000",
                     28275 => "01011001",
                     28276 => "01011010",
                     28277 => "01011010",
                     28278 => "00001000",
                     28279 => "00001001",
                     28280 => "00101000",
                     28281 => "00101001",
                     28282 => "00101010",
                     28283 => "00101011",
                     28284 => "00001110",
                     28285 => "00001111",
                     28286 => "11111100",
                     28287 => "11111100",
                     28288 => "11111100",
                     28289 => "11111100",
                     28290 => "00110010",
                     28291 => "00110011",
                     28292 => "00110100",
                     28293 => "00110101",
                     28294 => "11111100",
                     28295 => "11111100",
                     28296 => "11111100",
                     28297 => "11111100",
                     28298 => "00110110",
                     28299 => "00110111",
                     28300 => "00111000",
                     28301 => "00111001",
                     28302 => "11111100",
                     28303 => "11111100",
                     28304 => "11111100",
                     28305 => "11111100",
                     28306 => "00111010",
                     28307 => "00110111",
                     28308 => "00111011",
                     28309 => "00111100",
                     28310 => "11111100",
                     28311 => "11111100",
                     28312 => "11111100",
                     28313 => "11111100",
                     28314 => "00111101",
                     28315 => "00111110",
                     28316 => "00111111",
                     28317 => "01000000",
                     28318 => "11111100",
                     28319 => "11111100",
                     28320 => "11111100",
                     28321 => "11111100",
                     28322 => "00110010",
                     28323 => "01000001",
                     28324 => "01000010",
                     28325 => "01000011",
                     28326 => "11111100",
                     28327 => "11111100",
                     28328 => "11111100",
                     28329 => "11111100",
                     28330 => "00110010",
                     28331 => "00110011",
                     28332 => "01000100",
                     28333 => "01000101",
                     28334 => "11111100",
                     28335 => "11111100",
                     28336 => "11111100",
                     28337 => "11111100",
                     28338 => "00110010",
                     28339 => "00110011",
                     28340 => "01000100",
                     28341 => "01000111",
                     28342 => "11111100",
                     28343 => "11111100",
                     28344 => "11111100",
                     28345 => "11111100",
                     28346 => "00110010",
                     28347 => "00110011",
                     28348 => "01001000",
                     28349 => "01001001",
                     28350 => "11111100",
                     28351 => "11111100",
                     28352 => "11111100",
                     28353 => "11111100",
                     28354 => "00110010",
                     28355 => "00110011",
                     28356 => "10010000",
                     28357 => "10010001",
                     28358 => "11111100",
                     28359 => "11111100",
                     28360 => "11111100",
                     28361 => "11111100",
                     28362 => "00111010",
                     28363 => "00110111",
                     28364 => "10010010",
                     28365 => "10010011",
                     28366 => "11111100",
                     28367 => "11111100",
                     28368 => "11111100",
                     28369 => "11111100",
                     28370 => "10011110",
                     28371 => "10011110",
                     28372 => "10011111",
                     28373 => "10011111",
                     28374 => "11111100",
                     28375 => "11111100",
                     28376 => "11111100",
                     28377 => "11111100",
                     28378 => "00111010",
                     28379 => "00110111",
                     28380 => "01001111",
                     28381 => "01001111",
                     28382 => "11111100",
                     28383 => "11111100",
                     28384 => "00000000",
                     28385 => "00000001",
                     28386 => "01001100",
                     28387 => "01001101",
                     28388 => "01001110",
                     28389 => "01001110",
                     28390 => "00000000",
                     28391 => "00000001",
                     28392 => "01001100",
                     28393 => "01001101",
                     28394 => "01001010",
                     28395 => "01001010",
                     28396 => "01001011",
                     28397 => "01001011",
                     28398 => "00110001",
                     28399 => "01000110",
                     28400 => "10101101",
                     28401 => "10011110",
                     28402 => "00000111",
                     28403 => "11110000",
                     28404 => "00000101",
                     28405 => "10100101",
                     28406 => "00001001",
                     28407 => "01001010",
                     28408 => "10110000",
                     28409 => "01000000",
                     28410 => "10100101",
                     28411 => "00001110",
                     28412 => "11001001",
                     28413 => "00001011",
                     28414 => "11110000",
                     28415 => "01000111",
                     28416 => "10101101",
                     28417 => "00001011",
                     28418 => "00000111",
                     28419 => "11010000",
                     28420 => "00111100",
                     28421 => "10101100",
                     28422 => "00000100",
                     28423 => "00000111",
                     28424 => "11110000",
                     28425 => "00110001",
                     28426 => "10100101",
                     28427 => "00011101",
                     28428 => "11001001",
                     28429 => "00000000",
                     28430 => "11110000",
                     28431 => "00101011",
                     28432 => "00100000",
                     28433 => "00111011",
                     28434 => "11101111",
                     28435 => "10100101",
                     28436 => "00001001",
                     28437 => "00101001",
                     28438 => "00000100",
                     28439 => "11010000",
                     28440 => "00100001",
                     28441 => "10101010",
                     28442 => "10101100",
                     28443 => "11100100",
                     28444 => "00000110",
                     28445 => "10100101",
                     28446 => "00110011",
                     28447 => "01001010",
                     28448 => "10110000",
                     28449 => "00000100",
                     28450 => "11001000",
                     28451 => "11001000",
                     28452 => "11001000",
                     28453 => "11001000",
                     28454 => "10101101",
                     28455 => "01010100",
                     28456 => "00000111",
                     28457 => "11110000",
                     28458 => "00001001",
                     28459 => "10111001",
                     28460 => "00011001",
                     28461 => "00000010",
                     28462 => "11001101",
                     28463 => "10111100",
                     28464 => "11101110",
                     28465 => "11110000",
                     28466 => "00000111",
                     28467 => "11101000",
                     28468 => "10111101",
                     28469 => "11101110",
                     28470 => "11101110",
                     28471 => "10011001",
                     28472 => "00011001",
                     28473 => "00000010",
                     28474 => "01100000",
                     28475 => "00100000",
                     28476 => "11110011",
                     28477 => "11101111",
                     28478 => "01001100",
                     28479 => "01001100",
                     28480 => "11101111",
                     28481 => "00100000",
                     28482 => "10110111",
                     28483 => "11110000",
                     28484 => "01001100",
                     28485 => "01001100",
                     28486 => "11101111",
                     28487 => "10100000",
                     28488 => "00001110",
                     28489 => "10111001",
                     28490 => "00001110",
                     28491 => "11101110",
                     28492 => "10001101",
                     28493 => "11010101",
                     28494 => "00000110",
                     28495 => "10101001",
                     28496 => "00000100",
                     28497 => "00100000",
                     28498 => "11000101",
                     28499 => "11101111",
                     28500 => "00100000",
                     28501 => "11110000",
                     28502 => "11110000",
                     28503 => "10101101",
                     28504 => "00010001",
                     28505 => "00000111",
                     28506 => "11110000",
                     28507 => "00100101",
                     28508 => "10100000",
                     28509 => "00000000",
                     28510 => "10101101",
                     28511 => "10000001",
                     28512 => "00000111",
                     28513 => "11001101",
                     28514 => "00010001",
                     28515 => "00000111",
                     28516 => "10001100",
                     28517 => "00010001",
                     28518 => "00000111",
                     28519 => "10110000",
                     28520 => "00011000",
                     28521 => "10001101",
                     28522 => "00010001",
                     28523 => "00000111",
                     28524 => "10100000",
                     28525 => "00000111",
                     28526 => "10111001",
                     28527 => "00001110",
                     28528 => "11101110",
                     28529 => "10001101",
                     28530 => "11010101",
                     28531 => "00000110",
                     28532 => "10100000",
                     28533 => "00000100",
                     28534 => "10100101",
                     28535 => "01010111",
                     28536 => "00000101",
                     28537 => "00001100",
                     28538 => "11110000",
                     28539 => "00000001",
                     28540 => "10001000",
                     28541 => "10011000",
                     28542 => "00100000",
                     28543 => "11000101",
                     28544 => "11101111",
                     28545 => "10101101",
                     28546 => "11010000",
                     28547 => "00000011",
                     28548 => "01001010",
                     28549 => "01001010",
                     28550 => "01001010",
                     28551 => "01001010",
                     28552 => "10000101",
                     28553 => "00000000",
                     28554 => "10100010",
                     28555 => "00000011",
                     28556 => "10101101",
                     28557 => "11100100",
                     28558 => "00000110",
                     28559 => "00011000",
                     28560 => "01101001",
                     28561 => "00011000",
                     28562 => "10101000",
                     28563 => "10101001",
                     28564 => "11111000",
                     28565 => "01000110",
                     28566 => "00000000",
                     28567 => "10010000",
                     28568 => "00000011",
                     28569 => "00100000",
                     28570 => "11001000",
                     28571 => "11100101",
                     28572 => "10011000",
                     28573 => "00111000",
                     28574 => "11101001",
                     28575 => "00001000",
                     28576 => "10101000",
                     28577 => "11001010",
                     28578 => "00010000",
                     28579 => "11101111",
                     28580 => "01100000",
                     28581 => "01011000",
                     28582 => "00000001",
                     28583 => "00000000",
                     28584 => "01100000",
                     28585 => "11111111",
                     28586 => "00000100",
                     28587 => "10100010",
                     28588 => "00000101",
                     28589 => "10111101",
                     28590 => "10100101",
                     28591 => "11101111",
                     28592 => "10010101",
                     28593 => "00000010",
                     28594 => "11001010",
                     28595 => "00010000",
                     28596 => "11111000",
                     28597 => "10100010",
                     28598 => "10111000",
                     28599 => "10100000",
                     28600 => "00000100",
                     28601 => "00100000",
                     28602 => "11100011",
                     28603 => "11101111",
                     28604 => "10101101",
                     28605 => "00100110",
                     28606 => "00000010",
                     28607 => "00001001",
                     28608 => "01000000",
                     28609 => "10001101",
                     28610 => "00100010",
                     28611 => "00000010",
                     28612 => "01100000",
                     28613 => "10000101",
                     28614 => "00000111",
                     28615 => "10101101",
                     28616 => "10101101",
                     28617 => "00000011",
                     28618 => "10001101",
                     28619 => "01010101",
                     28620 => "00000111",
                     28621 => "10000101",
                     28622 => "00000101",
                     28623 => "10101101",
                     28624 => "10111000",
                     28625 => "00000011",
                     28626 => "10000101",
                     28627 => "00000010",
                     28628 => "10100101",
                     28629 => "00110011",
                     28630 => "10000101",
                     28631 => "00000011",
                     28632 => "10101101",
                     28633 => "11000100",
                     28634 => "00000011",
                     28635 => "10000101",
                     28636 => "00000100",
                     28637 => "10101110",
                     28638 => "11010101",
                     28639 => "00000110",
                     28640 => "10101100",
                     28641 => "11100100",
                     28642 => "00000110",
                     28643 => "10111101",
                     28644 => "00011110",
                     28645 => "11101110",
                     28646 => "10000101",
                     28647 => "00000000",
                     28648 => "10111101",
                     28649 => "00011111",
                     28650 => "11101110",
                     28651 => "00100000",
                     28652 => "10111001",
                     28653 => "11101011",
                     28654 => "11000110",
                     28655 => "00000111",
                     28656 => "11010000",
                     28657 => "11110001",
                     28658 => "01100000",
                     28659 => "10100101",
                     28660 => "00011101",
                     28661 => "11001001",
                     28662 => "00000011",
                     28663 => "11110000",
                     28664 => "01010010",
                     28665 => "11001001",
                     28666 => "00000010",
                     28667 => "11110000",
                     28668 => "00111110",
                     28669 => "11001001",
                     28670 => "00000001",
                     28671 => "11010000",
                     28672 => "00010001",
                     28673 => "10101101",
                     28674 => "00000100",
                     28675 => "00000111",
                     28676 => "11010000",
                     28677 => "01010001",
                     28678 => "10100000",
                     28679 => "00000110",
                     28680 => "10101101",
                     28681 => "00010100",
                     28682 => "00000111",
                     28683 => "11010000",
                     28684 => "00100010",
                     28685 => "10100000",
                     28686 => "00000000",
                     28687 => "01001100",
                     28688 => "00101111",
                     28689 => "11110000",
                     28690 => "10100000",
                     28691 => "00000110",
                     28692 => "10101101",
                     28693 => "00010100",
                     28694 => "00000111",
                     28695 => "11010000",
                     28696 => "00010110",
                     28697 => "10100000",
                     28698 => "00000010",
                     28699 => "10100101",
                     28700 => "01010111",
                     28701 => "00000101",
                     28702 => "00001100",
                     28703 => "11110000",
                     28704 => "00001110",
                     28705 => "10101101",
                     28706 => "00000000",
                     28707 => "00000111",
                     28708 => "11001001",
                     28709 => "00001010",
                     28710 => "10010000",
                     28711 => "00011011",
                     28712 => "10100101",
                     28713 => "01000101",
                     28714 => "00100101",
                     28715 => "00110011",
                     28716 => "11010000",
                     28717 => "00010101",
                     28718 => "11001000",
                     28719 => "00100000",
                     28720 => "10011000",
                     28721 => "11110000",
                     28722 => "10101001",
                     28723 => "00000000",
                     28724 => "10001101",
                     28725 => "00001101",
                     28726 => "00000111",
                     28727 => "10111001",
                     28728 => "00001110",
                     28729 => "11101110",
                     28730 => "01100000",
                     28731 => "10100000",
                     28732 => "00000100",
                     28733 => "00100000",
                     28734 => "10011000",
                     28735 => "11110000",
                     28736 => "01001100",
                     28737 => "01101001",
                     28738 => "11110000",
                     28739 => "10100000",
                     28740 => "00000100",
                     28741 => "00100000",
                     28742 => "10011000",
                     28743 => "11110000",
                     28744 => "01001100",
                     28745 => "01101111",
                     28746 => "11110000",
                     28747 => "10100000",
                     28748 => "00000101",
                     28749 => "10100101",
                     28750 => "10011111",
                     28751 => "11110000",
                     28752 => "11011110",
                     28753 => "00100000",
                     28754 => "10011000",
                     28755 => "11110000",
                     28756 => "01001100",
                     28757 => "01110100",
                     28758 => "11110000",
                     28759 => "10100000",
                     28760 => "00000001",
                     28761 => "00100000",
                     28762 => "10011000",
                     28763 => "11110000",
                     28764 => "10101101",
                     28765 => "10000010",
                     28766 => "00000111",
                     28767 => "00001101",
                     28768 => "00001101",
                     28769 => "00000111",
                     28770 => "11010000",
                     28771 => "00001011",
                     28772 => "10100101",
                     28773 => "00001010",
                     28774 => "00001010",
                     28775 => "10110000",
                     28776 => "00000110",
                     28777 => "10101101",
                     28778 => "00001101",
                     28779 => "00000111",
                     28780 => "01001100",
                     28781 => "11010111",
                     28782 => "11110000",
                     28783 => "10101001",
                     28784 => "00000011",
                     28785 => "01001100",
                     28786 => "01110110",
                     28787 => "11110000",
                     28788 => "10101001",
                     28789 => "00000010",
                     28790 => "10000101",
                     28791 => "00000000",
                     28792 => "00100000",
                     28793 => "01101001",
                     28794 => "11110000",
                     28795 => "01001000",
                     28796 => "10101101",
                     28797 => "10000001",
                     28798 => "00000111",
                     28799 => "11010000",
                     28800 => "00010101",
                     28801 => "10101101",
                     28802 => "00001100",
                     28803 => "00000111",
                     28804 => "10001101",
                     28805 => "10000001",
                     28806 => "00000111",
                     28807 => "10101101",
                     28808 => "00001101",
                     28809 => "00000111",
                     28810 => "00011000",
                     28811 => "01101001",
                     28812 => "00000001",
                     28813 => "11000101",
                     28814 => "00000000",
                     28815 => "10010000",
                     28816 => "00000010",
                     28817 => "10101001",
                     28818 => "00000000",
                     28819 => "10001101",
                     28820 => "00001101",
                     28821 => "00000111",
                     28822 => "01101000",
                     28823 => "01100000",
                     28824 => "10101101",
                     28825 => "01010100",
                     28826 => "00000111",
                     28827 => "11110000",
                     28828 => "00000101",
                     28829 => "10011000",
                     28830 => "00011000",
                     28831 => "01101001",
                     28832 => "00001000",
                     28833 => "10101000",
                     28834 => "01100000",
                     28835 => "00000000",
                     28836 => "00000001",
                     28837 => "00000000",
                     28838 => "00000001",
                     28839 => "00000000",
                     28840 => "00000001",
                     28841 => "00000010",
                     28842 => "00000000",
                     28843 => "00000001",
                     28844 => "00000010",
                     28845 => "00000010",
                     28846 => "00000000",
                     28847 => "00000010",
                     28848 => "00000000",
                     28849 => "00000010",
                     28850 => "00000000",
                     28851 => "00000010",
                     28852 => "00000000",
                     28853 => "00000010",
                     28854 => "00000000",
                     28855 => "10101100",
                     28856 => "00001101",
                     28857 => "00000111",
                     28858 => "10100101",
                     28859 => "00001001",
                     28860 => "00101001",
                     28861 => "00000011",
                     28862 => "11010000",
                     28863 => "00001101",
                     28864 => "11001000",
                     28865 => "11000000",
                     28866 => "00001010",
                     28867 => "10010000",
                     28868 => "00000101",
                     28869 => "10100000",
                     28870 => "00000000",
                     28871 => "10001100",
                     28872 => "00001011",
                     28873 => "00000111",
                     28874 => "10001100",
                     28875 => "00001101",
                     28876 => "00000111",
                     28877 => "10101101",
                     28878 => "01010100",
                     28879 => "00000111",
                     28880 => "11010000",
                     28881 => "00001100",
                     28882 => "10111001",
                     28883 => "10100011",
                     28884 => "11110000",
                     28885 => "10100000",
                     28886 => "00001111",
                     28887 => "00001010",
                     28888 => "00001010",
                     28889 => "00001010",
                     28890 => "01111001",
                     28891 => "00001110",
                     28892 => "11101110",
                     28893 => "01100000",
                     28894 => "10011000",
                     28895 => "00011000",
                     28896 => "01101001",
                     28897 => "00001010",
                     28898 => "10101010",
                     28899 => "10100000",
                     28900 => "00001001",
                     28901 => "10111101",
                     28902 => "10100011",
                     28903 => "11110000",
                     28904 => "11010000",
                     28905 => "00000010",
                     28906 => "10100000",
                     28907 => "00000001",
                     28908 => "10111001",
                     28909 => "00001110",
                     28910 => "11101110",
                     28911 => "01100000",
                     28912 => "10101100",
                     28913 => "11100100",
                     28914 => "00000110",
                     28915 => "10100101",
                     28916 => "00001110",
                     28917 => "11001001",
                     28918 => "00001011",
                     28919 => "11110000",
                     28920 => "00010011",
                     28921 => "10101101",
                     28922 => "11010101",
                     28923 => "00000110",
                     28924 => "11001001",
                     28925 => "01010000",
                     28926 => "11110000",
                     28927 => "00011110",
                     28928 => "11001001",
                     28929 => "10111000",
                     28930 => "11110000",
                     28931 => "00011010",
                     28932 => "11001001",
                     28933 => "11000000",
                     28934 => "11110000",
                     28935 => "00010110",
                     28936 => "11001001",
                     28937 => "11001000",
                     28938 => "11010000",
                     28939 => "00100100",
                     28940 => "10111001",
                     28941 => "00010010",
                     28942 => "00000010",
                     28943 => "00101001",
                     28944 => "00111111",
                     28945 => "10011001",
                     28946 => "00010010",
                     28947 => "00000010",
                     28948 => "10111001",
                     28949 => "00010110",
                     28950 => "00000010",
                     28951 => "00101001",
                     28952 => "00111111",
                     28953 => "00001001",
                     28954 => "01000000",
                     28955 => "10011001",
                     28956 => "00010110",
                     28957 => "00000010",
                     28958 => "10111001",
                     28959 => "00011010",
                     28960 => "00000010",
                     28961 => "00101001",
                     28962 => "00111111",
                     28963 => "10011001",
                     28964 => "00011010",
                     28965 => "00000010",
                     28966 => "10111001",
                     28967 => "00011110",
                     28968 => "00000010",
                     28969 => "00101001",
                     28970 => "00111111",
                     28971 => "00001001",
                     28972 => "01000000",
                     28973 => "10011001",
                     28974 => "00011110",
                     28975 => "00000010",
                     28976 => "01100000",
                     28977 => "10100010",
                     28978 => "00000000",
                     28979 => "10100000",
                     28980 => "00000000",
                     28981 => "01001100",
                     28982 => "01001001",
                     28983 => "11110001",
                     28984 => "10100000",
                     28985 => "00000001",
                     28986 => "00100000",
                     28987 => "10101111",
                     28988 => "11110001",
                     28989 => "10100000",
                     28990 => "00000011",
                     28991 => "01001100",
                     28992 => "01001001",
                     28993 => "11110001",
                     28994 => "10100000",
                     28995 => "00000000",
                     28996 => "00100000",
                     28997 => "10101111",
                     28998 => "11110001",
                     28999 => "10100000",
                     29000 => "00000010",
                     29001 => "00100000",
                     29002 => "01111000",
                     29003 => "11110001",
                     29004 => "10100110",
                     29005 => "00001000",
                     29006 => "01100000",
                     29007 => "10100000",
                     29008 => "00000010",
                     29009 => "00100000",
                     29010 => "10101111",
                     29011 => "11110001",
                     29012 => "10100000",
                     29013 => "00000110",
                     29014 => "01001100",
                     29015 => "01001001",
                     29016 => "11110001",
                     29017 => "10101001",
                     29018 => "00000001",
                     29019 => "10100000",
                     29020 => "00000001",
                     29021 => "01001100",
                     29022 => "01101100",
                     29023 => "11110001",
                     29024 => "10101001",
                     29025 => "00001001",
                     29026 => "10100000",
                     29027 => "00000100",
                     29028 => "00100000",
                     29029 => "01101100",
                     29030 => "11110001",
                     29031 => "11101000",
                     29032 => "11101000",
                     29033 => "10101001",
                     29034 => "00001001",
                     29035 => "11001000",
                     29036 => "10000110",
                     29037 => "00000000",
                     29038 => "00011000",
                     29039 => "01100101",
                     29040 => "00000000",
                     29041 => "10101010",
                     29042 => "00100000",
                     29043 => "01111000",
                     29044 => "11110001",
                     29045 => "10100110",
                     29046 => "00001000",
                     29047 => "01100000",
                     29048 => "10110101",
                     29049 => "11001110",
                     29050 => "10011001",
                     29051 => "10111000",
                     29052 => "00000011",
                     29053 => "10110101",
                     29054 => "10000110",
                     29055 => "00111000",
                     29056 => "11101101",
                     29057 => "00011100",
                     29058 => "00000111",
                     29059 => "10011001",
                     29060 => "10101101",
                     29061 => "00000011",
                     29062 => "01100000",
                     29063 => "10100010",
                     29064 => "00000000",
                     29065 => "10100000",
                     29066 => "00000000",
                     29067 => "01001100",
                     29068 => "11000111",
                     29069 => "11110001",
                     29070 => "10100000",
                     29071 => "00000000",
                     29072 => "00100000",
                     29073 => "10101111",
                     29074 => "11110001",
                     29075 => "10100000",
                     29076 => "00000010",
                     29077 => "01001100",
                     29078 => "11000111",
                     29079 => "11110001",
                     29080 => "10100000",
                     29081 => "00000001",
                     29082 => "00100000",
                     29083 => "10101111",
                     29084 => "11110001",
                     29085 => "10100000",
                     29086 => "00000011",
                     29087 => "01001100",
                     29088 => "11000111",
                     29089 => "11110001",
                     29090 => "10100000",
                     29091 => "00000010",
                     29092 => "00100000",
                     29093 => "10101111",
                     29094 => "11110001",
                     29095 => "10100000",
                     29096 => "00000110",
                     29097 => "01001100",
                     29098 => "11000111",
                     29099 => "11110001",
                     29100 => "00000111",
                     29101 => "00010110",
                     29102 => "00001101",
                     29103 => "10001010",
                     29104 => "00011000",
                     29105 => "01111001",
                     29106 => "10101100",
                     29107 => "11110001",
                     29108 => "10101010",
                     29109 => "01100000",
                     29110 => "10101001",
                     29111 => "00000001",
                     29112 => "10100000",
                     29113 => "00000001",
                     29114 => "01001100",
                     29115 => "11000001",
                     29116 => "11110001",
                     29117 => "10101001",
                     29118 => "00001001",
                     29119 => "10100000",
                     29120 => "00000100",
                     29121 => "10000110",
                     29122 => "00000000",
                     29123 => "00011000",
                     29124 => "01100101",
                     29125 => "00000000",
                     29126 => "10101010",
                     29127 => "10011000",
                     29128 => "01001000",
                     29129 => "00100000",
                     29130 => "11011110",
                     29131 => "11110001",
                     29132 => "00001010",
                     29133 => "00001010",
                     29134 => "00001010",
                     29135 => "00001010",
                     29136 => "00000101",
                     29137 => "00000000",
                     29138 => "10000101",
                     29139 => "00000000",
                     29140 => "01101000",
                     29141 => "10101000",
                     29142 => "10100101",
                     29143 => "00000000",
                     29144 => "10011001",
                     29145 => "11010000",
                     29146 => "00000011",
                     29147 => "10100110",
                     29148 => "00001000",
                     29149 => "01100000",
                     29150 => "00100000",
                     29151 => "11111101",
                     29152 => "11110001",
                     29153 => "01001010",
                     29154 => "01001010",
                     29155 => "01001010",
                     29156 => "01001010",
                     29157 => "10000101",
                     29158 => "00000000",
                     29159 => "01001100",
                     29160 => "01000000",
                     29161 => "11110010",
                     29162 => "01111111",
                     29163 => "00111111",
                     29164 => "00011111",
                     29165 => "00001111",
                     29166 => "00000111",
                     29167 => "00000011",
                     29168 => "00000001",
                     29169 => "00000000",
                     29170 => "10000000",
                     29171 => "11000000",
                     29172 => "11100000",
                     29173 => "11110000",
                     29174 => "11111000",
                     29175 => "11111100",
                     29176 => "11111110",
                     29177 => "11111111",
                     29178 => "00000111",
                     29179 => "00001111",
                     29180 => "00000111",
                     29181 => "10000110",
                     29182 => "00000100",
                     29183 => "10100000",
                     29184 => "00000001",
                     29185 => "10111001",
                     29186 => "00011100",
                     29187 => "00000111",
                     29188 => "00111000",
                     29189 => "11110101",
                     29190 => "10000110",
                     29191 => "10000101",
                     29192 => "00000111",
                     29193 => "10111001",
                     29194 => "00011010",
                     29195 => "00000111",
                     29196 => "11110101",
                     29197 => "01101101",
                     29198 => "10111110",
                     29199 => "11111010",
                     29200 => "11110001",
                     29201 => "11001001",
                     29202 => "00000000",
                     29203 => "00110000",
                     29204 => "00010000",
                     29205 => "10111110",
                     29206 => "11111011",
                     29207 => "11110001",
                     29208 => "11001001",
                     29209 => "00000001",
                     29210 => "00010000",
                     29211 => "00001001",
                     29212 => "10101001",
                     29213 => "00111000",
                     29214 => "10000101",
                     29215 => "00000110",
                     29216 => "10101001",
                     29217 => "00001000",
                     29218 => "00100000",
                     29219 => "01110100",
                     29220 => "11110010",
                     29221 => "10111101",
                     29222 => "11101010",
                     29223 => "11110001",
                     29224 => "10100110",
                     29225 => "00000100",
                     29226 => "11001001",
                     29227 => "00000000",
                     29228 => "11010000",
                     29229 => "00000011",
                     29230 => "10001000",
                     29231 => "00010000",
                     29232 => "11010000",
                     29233 => "01100000",
                     29234 => "00000000",
                     29235 => "00001000",
                     29236 => "00001100",
                     29237 => "00001110",
                     29238 => "00001111",
                     29239 => "00000111",
                     29240 => "00000011",
                     29241 => "00000001",
                     29242 => "00000000",
                     29243 => "00000100",
                     29244 => "00000000",
                     29245 => "00000100",
                     29246 => "11111111",
                     29247 => "00000000",
                     29248 => "10000110",
                     29249 => "00000100",
                     29250 => "10100000",
                     29251 => "00000001",
                     29252 => "10111001",
                     29253 => "00111110",
                     29254 => "11110010",
                     29255 => "00111000",
                     29256 => "11110101",
                     29257 => "11001110",
                     29258 => "10000101",
                     29259 => "00000111",
                     29260 => "10101001",
                     29261 => "00000001",
                     29262 => "11110101",
                     29263 => "10110101",
                     29264 => "10111110",
                     29265 => "00111011",
                     29266 => "11110010",
                     29267 => "11001001",
                     29268 => "00000000",
                     29269 => "00110000",
                     29270 => "00010000",
                     29271 => "10111110",
                     29272 => "00111100",
                     29273 => "11110010",
                     29274 => "11001001",
                     29275 => "00000001",
                     29276 => "00010000",
                     29277 => "00001001",
                     29278 => "10101001",
                     29279 => "00100000",
                     29280 => "10000101",
                     29281 => "00000110",
                     29282 => "10101001",
                     29283 => "00000100",
                     29284 => "00100000",
                     29285 => "01110100",
                     29286 => "11110010",
                     29287 => "10111101",
                     29288 => "00110010",
                     29289 => "11110010",
                     29290 => "10100110",
                     29291 => "00000100",
                     29292 => "11001001",
                     29293 => "00000000",
                     29294 => "11010000",
                     29295 => "00000011",
                     29296 => "10001000",
                     29297 => "00010000",
                     29298 => "11010001",
                     29299 => "01100000",
                     29300 => "10000101",
                     29301 => "00000101",
                     29302 => "10100101",
                     29303 => "00000111",
                     29304 => "11000101",
                     29305 => "00000110",
                     29306 => "10110000",
                     29307 => "00001100",
                     29308 => "01001010",
                     29309 => "01001010",
                     29310 => "01001010",
                     29311 => "00101001",
                     29312 => "00000111",
                     29313 => "11000000",
                     29314 => "00000001",
                     29315 => "10110000",
                     29316 => "00000010",
                     29317 => "01100101",
                     29318 => "00000101",
                     29319 => "10101010",
                     29320 => "01100000",
                     29321 => "10100101",
                     29322 => "00000011",
                     29323 => "01001010",
                     29324 => "01001010",
                     29325 => "10100101",
                     29326 => "00000000",
                     29327 => "10010000",
                     29328 => "00001100",
                     29329 => "10011001",
                     29330 => "00000101",
                     29331 => "00000010",
                     29332 => "10100101",
                     29333 => "00000001",
                     29334 => "10011001",
                     29335 => "00000001",
                     29336 => "00000010",
                     29337 => "10101001",
                     29338 => "01000000",
                     29339 => "11010000",
                     29340 => "00001010",
                     29341 => "10011001",
                     29342 => "00000001",
                     29343 => "00000010",
                     29344 => "10100101",
                     29345 => "00000001",
                     29346 => "10011001",
                     29347 => "00000101",
                     29348 => "00000010",
                     29349 => "10101001",
                     29350 => "00000000",
                     29351 => "00000101",
                     29352 => "00000100",
                     29353 => "10011001",
                     29354 => "00000010",
                     29355 => "00000010",
                     29356 => "10011001",
                     29357 => "00000110",
                     29358 => "00000010",
                     29359 => "10100101",
                     29360 => "00000010",
                     29361 => "10011001",
                     29362 => "00000000",
                     29363 => "00000010",
                     29364 => "10011001",
                     29365 => "00000100",
                     29366 => "00000010",
                     29367 => "10100101",
                     29368 => "00000101",
                     29369 => "10011001",
                     29370 => "00000011",
                     29371 => "00000010",
                     29372 => "00011000",
                     29373 => "01101001",
                     29374 => "00001000",
                     29375 => "10011001",
                     29376 => "00000111",
                     29377 => "00000010",
                     29378 => "10100101",
                     29379 => "00000010",
                     29380 => "00011000",
                     29381 => "01101001",
                     29382 => "00001000",
                     29383 => "10000101",
                     29384 => "00000010",
                     29385 => "10011000",
                     29386 => "00011000",
                     29387 => "01101001",
                     29388 => "00001000",
                     29389 => "10101000",
                     29390 => "11101000",
                     29391 => "11101000",
                     29392 => "01100000",
                     29393 => "10101101",
                     29394 => "01110000",
                     29395 => "00000111",
                     29396 => "11010000",
                     29397 => "00000100",
                     29398 => "10001101",
                     29399 => "00010101",
                     29400 => "01000000",
                     29401 => "01100000",
                     29402 => "10101001",
                     29403 => "11111111",
                     29404 => "10001101",
                     29405 => "00010111",
                     29406 => "01000000",
                     29407 => "10101001",
                     29408 => "00001111",
                     29409 => "10001101",
                     29410 => "00010101",
                     29411 => "01000000",
                     29412 => "10101101",
                     29413 => "11000110",
                     29414 => "00000111",
                     29415 => "11010000",
                     29416 => "00000110",
                     29417 => "10100101",
                     29418 => "11111010",
                     29419 => "11001001",
                     29420 => "00000001",
                     29421 => "11010000",
                     29422 => "01011101",
                     29423 => "10101101",
                     29424 => "10110010",
                     29425 => "00000111",
                     29426 => "11010000",
                     29427 => "00100011",
                     29428 => "10100101",
                     29429 => "11111010",
                     29430 => "11110000",
                     29431 => "01100110",
                     29432 => "10001101",
                     29433 => "10110010",
                     29434 => "00000111",
                     29435 => "10001101",
                     29436 => "11000110",
                     29437 => "00000111",
                     29438 => "10101001",
                     29439 => "00000000",
                     29440 => "10001101",
                     29441 => "00010101",
                     29442 => "01000000",
                     29443 => "10000101",
                     29444 => "11110001",
                     29445 => "10000101",
                     29446 => "11110010",
                     29447 => "10000101",
                     29448 => "11110011",
                     29449 => "10101001",
                     29450 => "00001111",
                     29451 => "10001101",
                     29452 => "00010101",
                     29453 => "01000000",
                     29454 => "10101001",
                     29455 => "00101010",
                     29456 => "10001101",
                     29457 => "10111011",
                     29458 => "00000111",
                     29459 => "10101001",
                     29460 => "01000100",
                     29461 => "11010000",
                     29462 => "00010001",
                     29463 => "10101101",
                     29464 => "10111011",
                     29465 => "00000111",
                     29466 => "11001001",
                     29467 => "00100100",
                     29468 => "11110000",
                     29469 => "00001000",
                     29470 => "11001001",
                     29471 => "00011110",
                     29472 => "11110000",
                     29473 => "11110001",
                     29474 => "11001001",
                     29475 => "00011000",
                     29476 => "11010000",
                     29477 => "00001001",
                     29478 => "10101001",
                     29479 => "01100100",
                     29480 => "10100010",
                     29481 => "10000100",
                     29482 => "10100000",
                     29483 => "01111111",
                     29484 => "00100000",
                     29485 => "10001001",
                     29486 => "11110011",
                     29487 => "11001110",
                     29488 => "10111011",
                     29489 => "00000111",
                     29490 => "11010000",
                     29491 => "00101010",
                     29492 => "10101001",
                     29493 => "00000000",
                     29494 => "10001101",
                     29495 => "00010101",
                     29496 => "01000000",
                     29497 => "10101101",
                     29498 => "10110010",
                     29499 => "00000111",
                     29500 => "11001001",
                     29501 => "00000010",
                     29502 => "11010000",
                     29503 => "00000101",
                     29504 => "10101001",
                     29505 => "00000000",
                     29506 => "10001101",
                     29507 => "11000110",
                     29508 => "00000111",
                     29509 => "10101001",
                     29510 => "00000000",
                     29511 => "10001101",
                     29512 => "10110010",
                     29513 => "00000111",
                     29514 => "11110000",
                     29515 => "00010010",
                     29516 => "00100000",
                     29517 => "00011100",
                     29518 => "11110100",
                     29519 => "00100000",
                     29520 => "01111101",
                     29521 => "11110101",
                     29522 => "00100000",
                     29523 => "01101000",
                     29524 => "11110110",
                     29525 => "00100000",
                     29526 => "10010101",
                     29527 => "11110110",
                     29528 => "10101001",
                     29529 => "00000000",
                     29530 => "10000101",
                     29531 => "11111011",
                     29532 => "10000101",
                     29533 => "11111100",
                     29534 => "10101001",
                     29535 => "00000000",
                     29536 => "10000101",
                     29537 => "11111111",
                     29538 => "10000101",
                     29539 => "11111110",
                     29540 => "10000101",
                     29541 => "11111101",
                     29542 => "10000101",
                     29543 => "11111010",
                     29544 => "10101100",
                     29545 => "11000000",
                     29546 => "00000111",
                     29547 => "10100101",
                     29548 => "11110100",
                     29549 => "00101001",
                     29550 => "00000011",
                     29551 => "11110000",
                     29552 => "00000111",
                     29553 => "11101110",
                     29554 => "11000000",
                     29555 => "00000111",
                     29556 => "11000000",
                     29557 => "00110000",
                     29558 => "10010000",
                     29559 => "00000110",
                     29560 => "10011000",
                     29561 => "11110000",
                     29562 => "00000011",
                     29563 => "11001110",
                     29564 => "11000000",
                     29565 => "00000111",
                     29566 => "10001100",
                     29567 => "00010001",
                     29568 => "01000000",
                     29569 => "01100000",
                     29570 => "10001100",
                     29571 => "00000001",
                     29572 => "01000000",
                     29573 => "10001110",
                     29574 => "00000000",
                     29575 => "01000000",
                     29576 => "01100000",
                     29577 => "00100000",
                     29578 => "10000010",
                     29579 => "11110011",
                     29580 => "10100010",
                     29581 => "00000000",
                     29582 => "10101000",
                     29583 => "10111001",
                     29584 => "00000001",
                     29585 => "11111111",
                     29586 => "11110000",
                     29587 => "00001011",
                     29588 => "10011101",
                     29589 => "00000010",
                     29590 => "01000000",
                     29591 => "10111001",
                     29592 => "00000000",
                     29593 => "11111111",
                     29594 => "00001001",
                     29595 => "00001000",
                     29596 => "10011101",
                     29597 => "00000011",
                     29598 => "01000000",
                     29599 => "01100000",
                     29600 => "10001110",
                     29601 => "00000100",
                     29602 => "01000000",
                     29603 => "10001100",
                     29604 => "00000101",
                     29605 => "01000000",
                     29606 => "01100000",
                     29607 => "00100000",
                     29608 => "10100000",
                     29609 => "11110011",
                     29610 => "10100010",
                     29611 => "00000100",
                     29612 => "11010000",
                     29613 => "11100000",
                     29614 => "10100010",
                     29615 => "00001000",
                     29616 => "11010000",
                     29617 => "11011100",
                     29618 => "10011111",
                     29619 => "10011011",
                     29620 => "10011000",
                     29621 => "10010110",
                     29622 => "10010101",
                     29623 => "10010100",
                     29624 => "10010010",
                     29625 => "10010000",
                     29626 => "10010000",
                     29627 => "10011010",
                     29628 => "10010111",
                     29629 => "10010101",
                     29630 => "10010011",
                     29631 => "10010010",
                     29632 => "10101001",
                     29633 => "01000000",
                     29634 => "10001101",
                     29635 => "10111011",
                     29636 => "00000111",
                     29637 => "10101001",
                     29638 => "01100010",
                     29639 => "00100000",
                     29640 => "10001100",
                     29641 => "11110011",
                     29642 => "10100010",
                     29643 => "10011001",
                     29644 => "11010000",
                     29645 => "00100101",
                     29646 => "10101001",
                     29647 => "00100110",
                     29648 => "11010000",
                     29649 => "00000010",
                     29650 => "10101001",
                     29651 => "00011000",
                     29652 => "10100010",
                     29653 => "10000010",
                     29654 => "10100000",
                     29655 => "10100111",
                     29656 => "00100000",
                     29657 => "10001001",
                     29658 => "11110011",
                     29659 => "10101001",
                     29660 => "00101000",
                     29661 => "10001101",
                     29662 => "10111011",
                     29663 => "00000111",
                     29664 => "10101101",
                     29665 => "10111011",
                     29666 => "00000111",
                     29667 => "11001001",
                     29668 => "00100101",
                     29669 => "11010000",
                     29670 => "00000110",
                     29671 => "10100010",
                     29672 => "01011111",
                     29673 => "10100000",
                     29674 => "11110110",
                     29675 => "11010000",
                     29676 => "00001000",
                     29677 => "11001001",
                     29678 => "00100000",
                     29679 => "11010000",
                     29680 => "00101001",
                     29681 => "10100010",
                     29682 => "01001000",
                     29683 => "10100000",
                     29684 => "10111100",
                     29685 => "00100000",
                     29686 => "10000010",
                     29687 => "11110011",
                     29688 => "11010000",
                     29689 => "00100000",
                     29690 => "10101001",
                     29691 => "00000101",
                     29692 => "10100000",
                     29693 => "10011001",
                     29694 => "11010000",
                     29695 => "00000100",
                     29696 => "10101001",
                     29697 => "00001010",
                     29698 => "10100000",
                     29699 => "10010011",
                     29700 => "10100010",
                     29701 => "10011110",
                     29702 => "10001101",
                     29703 => "10111011",
                     29704 => "00000111",
                     29705 => "10101001",
                     29706 => "00001100",
                     29707 => "00100000",
                     29708 => "10001001",
                     29709 => "11110011",
                     29710 => "10101101",
                     29711 => "10111011",
                     29712 => "00000111",
                     29713 => "11001001",
                     29714 => "00000110",
                     29715 => "11010000",
                     29716 => "00000101",
                     29717 => "10101001",
                     29718 => "10111011",
                     29719 => "10001101",
                     29720 => "00000001",
                     29721 => "01000000",
                     29722 => "11010000",
                     29723 => "01100000",
                     29724 => "10100100",
                     29725 => "11111111",
                     29726 => "11110000",
                     29727 => "00100000",
                     29728 => "10000100",
                     29729 => "11110001",
                     29730 => "00110000",
                     29731 => "10101010",
                     29732 => "01000110",
                     29733 => "11111111",
                     29734 => "10110000",
                     29735 => "10101010",
                     29736 => "01000110",
                     29737 => "11111111",
                     29738 => "10110000",
                     29739 => "11010100",
                     29740 => "01000110",
                     29741 => "11111111",
                     29742 => "10110000",
                     29743 => "00101100",
                     29744 => "01000110",
                     29745 => "11111111",
                     29746 => "10110000",
                     29747 => "01001010",
                     29748 => "01000110",
                     29749 => "11111111",
                     29750 => "10110000",
                     29751 => "01111111",
                     29752 => "01000110",
                     29753 => "11111111",
                     29754 => "10110000",
                     29755 => "10111110",
                     29756 => "01000110",
                     29757 => "11111111",
                     29758 => "10110000",
                     29759 => "10000000",
                     29760 => "10100101",
                     29761 => "11110001",
                     29762 => "11110000",
                     29763 => "00010111",
                     29764 => "00110000",
                     29765 => "10011010",
                     29766 => "01001010",
                     29767 => "10110000",
                     29768 => "10010111",
                     29769 => "01001010",
                     29770 => "10110000",
                     29771 => "11000010",
                     29772 => "01001010",
                     29773 => "10110000",
                     29774 => "00011011",
                     29775 => "01001010",
                     29776 => "10110000",
                     29777 => "00111100",
                     29778 => "01001010",
                     29779 => "10110000",
                     29780 => "01100111",
                     29781 => "01001010",
                     29782 => "10110000",
                     29783 => "10110110",
                     29784 => "01001010",
                     29785 => "10110000",
                     29786 => "01001000",
                     29787 => "01100000",
                     29788 => "10101001",
                     29789 => "00001110",
                     29790 => "10001101",
                     29791 => "10111011",
                     29792 => "00000111",
                     29793 => "10100000",
                     29794 => "10011100",
                     29795 => "10100010",
                     29796 => "10011110",
                     29797 => "10101001",
                     29798 => "00100110",
                     29799 => "00100000",
                     29800 => "10001001",
                     29801 => "11110011",
                     29802 => "10101100",
                     29803 => "10111011",
                     29804 => "00000111",
                     29805 => "10111001",
                     29806 => "10110001",
                     29807 => "11110011",
                     29808 => "10001101",
                     29809 => "00000000",
                     29810 => "01000000",
                     29811 => "11000000",
                     29812 => "00000110",
                     29813 => "11010000",
                     29814 => "00000101",
                     29815 => "10101001",
                     29816 => "10011110",
                     29817 => "10001101",
                     29818 => "00000010",
                     29819 => "01000000",
                     29820 => "11010000",
                     29821 => "00100101",
                     29822 => "10101001",
                     29823 => "00001110",
                     29824 => "10100000",
                     29825 => "11001011",
                     29826 => "10100010",
                     29827 => "10011111",
                     29828 => "10001101",
                     29829 => "10111011",
                     29830 => "00000111",
                     29831 => "10101001",
                     29832 => "00101000",
                     29833 => "00100000",
                     29834 => "10001001",
                     29835 => "11110011",
                     29836 => "11010000",
                     29837 => "00010101",
                     29838 => "10101100",
                     29839 => "10111011",
                     29840 => "00000111",
                     29841 => "11000000",
                     29842 => "00001000",
                     29843 => "11010000",
                     29844 => "00001001",
                     29845 => "10101001",
                     29846 => "10100000",
                     29847 => "10001101",
                     29848 => "00000010",
                     29849 => "01000000",
                     29850 => "10101001",
                     29851 => "10011111",
                     29852 => "11010000",
                     29853 => "00000010",
                     29854 => "10101001",
                     29855 => "10010000",
                     29856 => "10001101",
                     29857 => "00000000",
                     29858 => "01000000",
                     29859 => "11001110",
                     29860 => "10111011",
                     29861 => "00000111",
                     29862 => "11010000",
                     29863 => "00001110",
                     29864 => "10100010",
                     29865 => "00000000",
                     29866 => "10000110",
                     29867 => "11110001",
                     29868 => "10100010",
                     29869 => "00001110",
                     29870 => "10001110",
                     29871 => "00010101",
                     29872 => "01000000",
                     29873 => "10100010",
                     29874 => "00001111",
                     29875 => "10001110",
                     29876 => "00010101",
                     29877 => "01000000",
                     29878 => "01100000",
                     29879 => "10101001",
                     29880 => "00101111",
                     29881 => "10001101",
                     29882 => "10111011",
                     29883 => "00000111",
                     29884 => "10101101",
                     29885 => "10111011",
                     29886 => "00000111",
                     29887 => "01001010",
                     29888 => "10110000",
                     29889 => "00010000",
                     29890 => "01001010",
                     29891 => "10110000",
                     29892 => "00001101",
                     29893 => "00101001",
                     29894 => "00000010",
                     29895 => "11110000",
                     29896 => "00001001",
                     29897 => "10100000",
                     29898 => "10010001",
                     29899 => "10100010",
                     29900 => "10011010",
                     29901 => "10101001",
                     29902 => "01000100",
                     29903 => "00100000",
                     29904 => "10001001",
                     29905 => "11110011",
                     29906 => "01001100",
                     29907 => "10100011",
                     29908 => "11110100",
                     29909 => "01011000",
                     29910 => "00000010",
                     29911 => "01010100",
                     29912 => "01010110",
                     29913 => "01001110",
                     29914 => "01000100",
                     29915 => "01001100",
                     29916 => "01010010",
                     29917 => "01001100",
                     29918 => "01001000",
                     29919 => "00111110",
                     29920 => "00110110",
                     29921 => "00111110",
                     29922 => "00110110",
                     29923 => "00110000",
                     29924 => "00101000",
                     29925 => "01001010",
                     29926 => "01010000",
                     29927 => "01001010",
                     29928 => "01100100",
                     29929 => "00111100",
                     29930 => "00110010",
                     29931 => "00111100",
                     29932 => "00110010",
                     29933 => "00101100",
                     29934 => "00100100",
                     29935 => "00111010",
                     29936 => "01100100",
                     29937 => "00111010",
                     29938 => "00110100",
                     29939 => "00101100",
                     29940 => "00100010",
                     29941 => "00101100",
                     29942 => "00100010",
                     29943 => "00011100",
                     29944 => "00010100",
                     29945 => "00010100",
                     29946 => "00000100",
                     29947 => "00100010",
                     29948 => "00100100",
                     29949 => "00010110",
                     29950 => "00000100",
                     29951 => "00100100",
                     29952 => "00100110",
                     29953 => "00011000",
                     29954 => "00000100",
                     29955 => "00100110",
                     29956 => "00101000",
                     29957 => "00011010",
                     29958 => "00000100",
                     29959 => "00101000",
                     29960 => "00101010",
                     29961 => "00011100",
                     29962 => "00000100",
                     29963 => "00101010",
                     29964 => "00101100",
                     29965 => "00011110",
                     29966 => "00000100",
                     29967 => "00101100",
                     29968 => "00101110",
                     29969 => "00100000",
                     29970 => "00000100",
                     29971 => "00101110",
                     29972 => "00110000",
                     29973 => "00100010",
                     29974 => "00000100",
                     29975 => "00110000",
                     29976 => "00110010",
                     29977 => "10101001",
                     29978 => "00110101",
                     29979 => "10100010",
                     29980 => "10001101",
                     29981 => "11010000",
                     29982 => "00000100",
                     29983 => "10101001",
                     29984 => "00000110",
                     29985 => "10100010",
                     29986 => "10011000",
                     29987 => "10001101",
                     29988 => "10111101",
                     29989 => "00000111",
                     29990 => "10100000",
                     29991 => "01111111",
                     29992 => "10101001",
                     29993 => "01000010",
                     29994 => "00100000",
                     29995 => "10100111",
                     29996 => "11110011",
                     29997 => "10101101",
                     29998 => "10111101",
                     29999 => "00000111",
                     30000 => "11001001",
                     30001 => "00110000",
                     30002 => "11010000",
                     30003 => "00000101",
                     30004 => "10101001",
                     30005 => "01001110",
                     30006 => "10001101",
                     30007 => "00000110",
                     30008 => "01000000",
                     30009 => "11010000",
                     30010 => "00101110",
                     30011 => "10101001",
                     30012 => "00100000",
                     30013 => "10001101",
                     30014 => "10111101",
                     30015 => "00000111",
                     30016 => "10100000",
                     30017 => "10010100",
                     30018 => "10101001",
                     30019 => "01011110",
                     30020 => "11010000",
                     30021 => "00001011",
                     30022 => "10101101",
                     30023 => "10111101",
                     30024 => "00000111",
                     30025 => "11001001",
                     30026 => "00011000",
                     30027 => "11010000",
                     30028 => "00011100",
                     30029 => "10100000",
                     30030 => "10010011",
                     30031 => "10101001",
                     30032 => "00011000",
                     30033 => "11010000",
                     30034 => "01111111",
                     30035 => "10101001",
                     30036 => "00110110",
                     30037 => "10001101",
                     30038 => "10111101",
                     30039 => "00000111",
                     30040 => "10101101",
                     30041 => "10111101",
                     30042 => "00000111",
                     30043 => "01001010",
                     30044 => "10110000",
                     30045 => "00001011",
                     30046 => "10101000",
                     30047 => "10111001",
                     30048 => "11011010",
                     30049 => "11110100",
                     30050 => "10100010",
                     30051 => "01011101",
                     30052 => "10100000",
                     30053 => "01111111",
                     30054 => "00100000",
                     30055 => "10100111",
                     30056 => "11110011",
                     30057 => "11001110",
                     30058 => "10111101",
                     30059 => "00000111",
                     30060 => "11010000",
                     30061 => "00001110",
                     30062 => "10100010",
                     30063 => "00000000",
                     30064 => "10000110",
                     30065 => "11110010",
                     30066 => "10100010",
                     30067 => "00001101",
                     30068 => "10001110",
                     30069 => "00010101",
                     30070 => "01000000",
                     30071 => "10100010",
                     30072 => "00001111",
                     30073 => "10001110",
                     30074 => "00010101",
                     30075 => "01000000",
                     30076 => "01100000",
                     30077 => "10100101",
                     30078 => "11110010",
                     30079 => "00101001",
                     30080 => "01000000",
                     30081 => "11010000",
                     30082 => "01100101",
                     30083 => "10100100",
                     30084 => "11111110",
                     30085 => "11110000",
                     30086 => "00100000",
                     30087 => "10000100",
                     30088 => "11110010",
                     30089 => "00110000",
                     30090 => "00111110",
                     30091 => "01000110",
                     30092 => "11111110",
                     30093 => "10110000",
                     30094 => "10001010",
                     30095 => "01000110",
                     30096 => "11111110",
                     30097 => "10110000",
                     30098 => "01101010",
                     30099 => "01000110",
                     30100 => "11111110",
                     30101 => "10110000",
                     30102 => "01101010",
                     30103 => "01000110",
                     30104 => "11111110",
                     30105 => "10110000",
                     30106 => "10100000",
                     30107 => "01000110",
                     30108 => "11111110",
                     30109 => "10110000",
                     30110 => "10000000",
                     30111 => "01000110",
                     30112 => "11111110",
                     30113 => "10110000",
                     30114 => "10110000",
                     30115 => "01000110",
                     30116 => "11111110",
                     30117 => "10110000",
                     30118 => "00111100",
                     30119 => "10100101",
                     30120 => "11110010",
                     30121 => "11110000",
                     30122 => "00010111",
                     30123 => "00110000",
                     30124 => "00100111",
                     30125 => "01001010",
                     30126 => "10110000",
                     30127 => "00010011",
                     30128 => "01001010",
                     30129 => "10110000",
                     30130 => "01011101",
                     30131 => "01001010",
                     30132 => "10110000",
                     30133 => "01011010",
                     30134 => "01001010",
                     30135 => "10110000",
                     30136 => "10001101",
                     30137 => "01001010",
                     30138 => "10110000",
                     30139 => "00000111",
                     30140 => "01001010",
                     30141 => "10110000",
                     30142 => "10011001",
                     30143 => "01001010",
                     30144 => "10110000",
                     30145 => "00100110",
                     30146 => "01100000",
                     30147 => "01001100",
                     30148 => "00101101",
                     30149 => "11110101",
                     30150 => "01001100",
                     30151 => "01101001",
                     30152 => "11110101",
                     30153 => "10101001",
                     30154 => "00111000",
                     30155 => "10001101",
                     30156 => "10111101",
                     30157 => "00000111",
                     30158 => "10100000",
                     30159 => "11000100",
                     30160 => "10101001",
                     30161 => "00011000",
                     30162 => "11010000",
                     30163 => "00001011",
                     30164 => "10101101",
                     30165 => "10111101",
                     30166 => "00000111",
                     30167 => "11001001",
                     30168 => "00001000",
                     30169 => "11010000",
                     30170 => "10001110",
                     30171 => "10100000",
                     30172 => "10100100",
                     30173 => "10101001",
                     30174 => "01011010",
                     30175 => "10100010",
                     30176 => "10011111",
                     30177 => "11010000",
                     30178 => "10000011",
                     30179 => "10101001",
                     30180 => "00110000",
                     30181 => "10001101",
                     30182 => "10111101",
                     30183 => "00000111",
                     30184 => "10101101",
                     30185 => "10111101",
                     30186 => "00000111",
                     30187 => "10100010",
                     30188 => "00000011",
                     30189 => "01001010",
                     30190 => "10110000",
                     30191 => "11010110",
                     30192 => "11001010",
                     30193 => "11010000",
                     30194 => "11111010",
                     30195 => "10101000",
                     30196 => "10111001",
                     30197 => "11010100",
                     30198 => "11110100",
                     30199 => "10100010",
                     30200 => "10000010",
                     30201 => "10100000",
                     30202 => "01111111",
                     30203 => "11010000",
                     30204 => "11100100",
                     30205 => "10101001",
                     30206 => "00010000",
                     30207 => "11010000",
                     30208 => "00000010",
                     30209 => "10101001",
                     30210 => "00100000",
                     30211 => "10001101",
                     30212 => "10111101",
                     30213 => "00000111",
                     30214 => "10101001",
                     30215 => "01111111",
                     30216 => "10001101",
                     30217 => "00000101",
                     30218 => "01000000",
                     30219 => "10101001",
                     30220 => "00000000",
                     30221 => "10001101",
                     30222 => "10111110",
                     30223 => "00000111",
                     30224 => "11101110",
                     30225 => "10111110",
                     30226 => "00000111",
                     30227 => "10101101",
                     30228 => "10111110",
                     30229 => "00000111",
                     30230 => "01001010",
                     30231 => "10101000",
                     30232 => "11001100",
                     30233 => "10111101",
                     30234 => "00000111",
                     30235 => "11110000",
                     30236 => "00001100",
                     30237 => "10101001",
                     30238 => "10011101",
                     30239 => "10001101",
                     30240 => "00000100",
                     30241 => "01000000",
                     30242 => "10111001",
                     30243 => "11111001",
                     30244 => "11110100",
                     30245 => "00100000",
                     30246 => "10101010",
                     30247 => "11110011",
                     30248 => "01100000",
                     30249 => "01001100",
                     30250 => "01101110",
                     30251 => "11110101",
                     30252 => "00000001",
                     30253 => "00001110",
                     30254 => "00001110",
                     30255 => "00001101",
                     30256 => "00001011",
                     30257 => "00000110",
                     30258 => "00001100",
                     30259 => "00001111",
                     30260 => "00001010",
                     30261 => "00001001",
                     30262 => "00000011",
                     30263 => "00001101",
                     30264 => "00001000",
                     30265 => "00001101",
                     30266 => "00000110",
                     30267 => "00001100",
                     30268 => "10101001",
                     30269 => "00100000",
                     30270 => "10001101",
                     30271 => "10111111",
                     30272 => "00000111",
                     30273 => "10101101",
                     30274 => "10111111",
                     30275 => "00000111",
                     30276 => "01001010",
                     30277 => "10010000",
                     30278 => "00010010",
                     30279 => "10101000",
                     30280 => "10111110",
                     30281 => "00101100",
                     30282 => "11110110",
                     30283 => "10111001",
                     30284 => "11101010",
                     30285 => "11111111",
                     30286 => "10001101",
                     30287 => "00001100",
                     30288 => "01000000",
                     30289 => "10001110",
                     30290 => "00001110",
                     30291 => "01000000",
                     30292 => "10101001",
                     30293 => "00011000",
                     30294 => "10001101",
                     30295 => "00001111",
                     30296 => "01000000",
                     30297 => "11001110",
                     30298 => "10111111",
                     30299 => "00000111",
                     30300 => "11010000",
                     30301 => "00001001",
                     30302 => "10101001",
                     30303 => "11110000",
                     30304 => "10001101",
                     30305 => "00001100",
                     30306 => "01000000",
                     30307 => "10101001",
                     30308 => "00000000",
                     30309 => "10000101",
                     30310 => "11110011",
                     30311 => "01100000",
                     30312 => "10100100",
                     30313 => "11111101",
                     30314 => "11110000",
                     30315 => "00001010",
                     30316 => "10000100",
                     30317 => "11110011",
                     30318 => "01000110",
                     30319 => "11111101",
                     30320 => "10110000",
                     30321 => "11001010",
                     30322 => "01000110",
                     30323 => "11111101",
                     30324 => "10110000",
                     30325 => "00001011",
                     30326 => "10100101",
                     30327 => "11110011",
                     30328 => "11110000",
                     30329 => "00000110",
                     30330 => "01001010",
                     30331 => "10110000",
                     30332 => "11000100",
                     30333 => "01001010",
                     30334 => "10110000",
                     30335 => "00000110",
                     30336 => "01100000",
                     30337 => "10101001",
                     30338 => "01000000",
                     30339 => "10001101",
                     30340 => "10111111",
                     30341 => "00000111",
                     30342 => "10101101",
                     30343 => "10111111",
                     30344 => "00000111",
                     30345 => "01001010",
                     30346 => "10101000",
                     30347 => "10100010",
                     30348 => "00001111",
                     30349 => "10111001",
                     30350 => "11001001",
                     30351 => "11111111",
                     30352 => "11010000",
                     30353 => "10111100",
                     30354 => "01001100",
                     30355 => "00111011",
                     30356 => "11110111",
                     30357 => "10100101",
                     30358 => "11111100",
                     30359 => "11010000",
                     30360 => "00001100",
                     30361 => "10100101",
                     30362 => "11111011",
                     30363 => "11010000",
                     30364 => "00101100",
                     30365 => "10101101",
                     30366 => "10110001",
                     30367 => "00000111",
                     30368 => "00000101",
                     30369 => "11110100",
                     30370 => "11010000",
                     30371 => "11101110",
                     30372 => "01100000",
                     30373 => "10001101",
                     30374 => "10110001",
                     30375 => "00000111",
                     30376 => "11001001",
                     30377 => "00000001",
                     30378 => "11010000",
                     30379 => "00000110",
                     30380 => "00100000",
                     30381 => "10101000",
                     30382 => "11110100",
                     30383 => "00100000",
                     30384 => "01110010",
                     30385 => "11110101",
                     30386 => "10100110",
                     30387 => "11110100",
                     30388 => "10001110",
                     30389 => "11000101",
                     30390 => "00000111",
                     30391 => "10100000",
                     30392 => "00000000",
                     30393 => "10001100",
                     30394 => "11000100",
                     30395 => "00000111",
                     30396 => "10000100",
                     30397 => "11110100",
                     30398 => "11001001",
                     30399 => "01000000",
                     30400 => "11010000",
                     30401 => "00110000",
                     30402 => "10100010",
                     30403 => "00001000",
                     30404 => "10001110",
                     30405 => "11000100",
                     30406 => "00000111",
                     30407 => "11010000",
                     30408 => "00101001",
                     30409 => "11001001",
                     30410 => "00000100",
                     30411 => "11010000",
                     30412 => "00000011",
                     30413 => "00100000",
                     30414 => "10101000",
                     30415 => "11110100",
                     30416 => "10100000",
                     30417 => "00010000",
                     30418 => "10001100",
                     30419 => "11000111",
                     30420 => "00000111",
                     30421 => "10100000",
                     30422 => "00000000",
                     30423 => "10001100",
                     30424 => "10110001",
                     30425 => "00000111",
                     30426 => "10000101",
                     30427 => "11110100",
                     30428 => "11001001",
                     30429 => "00000001",
                     30430 => "11010000",
                     30431 => "00001110",
                     30432 => "11101110",
                     30433 => "11000111",
                     30434 => "00000111",
                     30435 => "10101100",
                     30436 => "11000111",
                     30437 => "00000111",
                     30438 => "11000000",
                     30439 => "00110010",
                     30440 => "11010000",
                     30441 => "00001100",
                     30442 => "10100000",
                     30443 => "00010001",
                     30444 => "11010000",
                     30445 => "11100100",
                     30446 => "10100000",
                     30447 => "00001000",
                     30448 => "10000100",
                     30449 => "11110111",
                     30450 => "11001000",
                     30451 => "01001010",
                     30452 => "10010000",
                     30453 => "11111100",
                     30454 => "10111001",
                     30455 => "00001101",
                     30456 => "11111001",
                     30457 => "10101000",
                     30458 => "10111001",
                     30459 => "00001110",
                     30460 => "11111001",
                     30461 => "10000101",
                     30462 => "11110000",
                     30463 => "10111001",
                     30464 => "00001111",
                     30465 => "11111001",
                     30466 => "10000101",
                     30467 => "11110101",
                     30468 => "10111001",
                     30469 => "00010000",
                     30470 => "11111001",
                     30471 => "10000101",
                     30472 => "11110110",
                     30473 => "10111001",
                     30474 => "00010001",
                     30475 => "11111001",
                     30476 => "10000101",
                     30477 => "11111001",
                     30478 => "10111001",
                     30479 => "00010010",
                     30480 => "11111001",
                     30481 => "10000101",
                     30482 => "11111000",
                     30483 => "10111001",
                     30484 => "00010011",
                     30485 => "11111001",
                     30486 => "10001101",
                     30487 => "10110000",
                     30488 => "00000111",
                     30489 => "10001101",
                     30490 => "11000001",
                     30491 => "00000111",
                     30492 => "10101001",
                     30493 => "00000001",
                     30494 => "10001101",
                     30495 => "10110100",
                     30496 => "00000111",
                     30497 => "10001101",
                     30498 => "10110110",
                     30499 => "00000111",
                     30500 => "10001101",
                     30501 => "10111001",
                     30502 => "00000111",
                     30503 => "10001101",
                     30504 => "10111010",
                     30505 => "00000111",
                     30506 => "10101001",
                     30507 => "00000000",
                     30508 => "10000101",
                     30509 => "11110111",
                     30510 => "10001101",
                     30511 => "11001010",
                     30512 => "00000111",
                     30513 => "10101001",
                     30514 => "00001011",
                     30515 => "10001101",
                     30516 => "00010101",
                     30517 => "01000000",
                     30518 => "10101001",
                     30519 => "00001111",
                     30520 => "10001101",
                     30521 => "00010101",
                     30522 => "01000000",
                     30523 => "11001110",
                     30524 => "10110100",
                     30525 => "00000111",
                     30526 => "11010000",
                     30527 => "01011111",
                     30528 => "10100100",
                     30529 => "11110111",
                     30530 => "11100110",
                     30531 => "11110111",
                     30532 => "10110001",
                     30533 => "11110101",
                     30534 => "11110000",
                     30535 => "00000100",
                     30536 => "00010000",
                     30537 => "00111101",
                     30538 => "11010000",
                     30539 => "00101111",
                     30540 => "10101101",
                     30541 => "10110001",
                     30542 => "00000111",
                     30543 => "11001001",
                     30544 => "01000000",
                     30545 => "11010000",
                     30546 => "00000101",
                     30547 => "10101101",
                     30548 => "11000101",
                     30549 => "00000111",
                     30550 => "11010000",
                     30551 => "00011101",
                     30552 => "00101001",
                     30553 => "00000100",
                     30554 => "11010000",
                     30555 => "00011100",
                     30556 => "10100101",
                     30557 => "11110100",
                     30558 => "00101001",
                     30559 => "01011111",
                     30560 => "11010000",
                     30561 => "00010011",
                     30562 => "10101001",
                     30563 => "00000000",
                     30564 => "10000101",
                     30565 => "11110100",
                     30566 => "10001101",
                     30567 => "10110001",
                     30568 => "00000111",
                     30569 => "10001101",
                     30570 => "00001000",
                     30571 => "01000000",
                     30572 => "10101001",
                     30573 => "10010000",
                     30574 => "10001101",
                     30575 => "00000000",
                     30576 => "01000000",
                     30577 => "10001101",
                     30578 => "00000100",
                     30579 => "01000000",
                     30580 => "01100000",
                     30581 => "01001100",
                     30582 => "11010101",
                     30583 => "11110110",
                     30584 => "01001100",
                     30585 => "10100101",
                     30586 => "11110110",
                     30587 => "00100000",
                     30588 => "11001100",
                     30589 => "11111000",
                     30590 => "10001101",
                     30591 => "10110011",
                     30592 => "00000111",
                     30593 => "10100100",
                     30594 => "11110111",
                     30595 => "11100110",
                     30596 => "11110111",
                     30597 => "10110001",
                     30598 => "11110101",
                     30599 => "10100110",
                     30600 => "11110010",
                     30601 => "11010000",
                     30602 => "00001110",
                     30603 => "00100000",
                     30604 => "10101010",
                     30605 => "11110011",
                     30606 => "11110000",
                     30607 => "00000011",
                     30608 => "00100000",
                     30609 => "11011001",
                     30610 => "11111000",
                     30611 => "10001101",
                     30612 => "10110101",
                     30613 => "00000111",
                     30614 => "00100000",
                     30615 => "10100000",
                     30616 => "11110011",
                     30617 => "10101101",
                     30618 => "10110011",
                     30619 => "00000111",
                     30620 => "10001101",
                     30621 => "10110100",
                     30622 => "00000111",
                     30623 => "10100101",
                     30624 => "11110010",
                     30625 => "11010000",
                     30626 => "00011010",
                     30627 => "10101101",
                     30628 => "10110001",
                     30629 => "00000111",
                     30630 => "00101001",
                     30631 => "10010001",
                     30632 => "11010000",
                     30633 => "00010011",
                     30634 => "10101100",
                     30635 => "10110101",
                     30636 => "00000111",
                     30637 => "11110000",
                     30638 => "00000011",
                     30639 => "11001110",
                     30640 => "10110101",
                     30641 => "00000111",
                     30642 => "00100000",
                     30643 => "11110101",
                     30644 => "11111000",
                     30645 => "10001101",
                     30646 => "00000100",
                     30647 => "01000000",
                     30648 => "10100010",
                     30649 => "01111111",
                     30650 => "10001110",
                     30651 => "00000101",
                     30652 => "01000000",
                     30653 => "10100100",
                     30654 => "11111000",
                     30655 => "11110000",
                     30656 => "01011010",
                     30657 => "11001110",
                     30658 => "10110110",
                     30659 => "00000111",
                     30660 => "11010000",
                     30661 => "00110010",
                     30662 => "10100100",
                     30663 => "11111000",
                     30664 => "11100110",
                     30665 => "11111000",
                     30666 => "10110001",
                     30667 => "11110101",
                     30668 => "11010000",
                     30669 => "00001111",
                     30670 => "10101001",
                     30671 => "10000011",
                     30672 => "10001101",
                     30673 => "00000000",
                     30674 => "01000000",
                     30675 => "10101001",
                     30676 => "10010100",
                     30677 => "10001101",
                     30678 => "00000001",
                     30679 => "01000000",
                     30680 => "10001101",
                     30681 => "11001010",
                     30682 => "00000111",
                     30683 => "11010000",
                     30684 => "11101001",
                     30685 => "00100000",
                     30686 => "11000110",
                     30687 => "11111000",
                     30688 => "10001101",
                     30689 => "10110110",
                     30690 => "00000111",
                     30691 => "10100100",
                     30692 => "11110001",
                     30693 => "11010000",
                     30694 => "00110100",
                     30695 => "10001010",
                     30696 => "00101001",
                     30697 => "00111110",
                     30698 => "00100000",
                     30699 => "10001100",
                     30700 => "11110011",
                     30701 => "11110000",
                     30702 => "00000011",
                     30703 => "00100000",
                     30704 => "11011001",
                     30705 => "11111000",
                     30706 => "10001101",
                     30707 => "10110111",
                     30708 => "00000111",
                     30709 => "00100000",
                     30710 => "10000010",
                     30711 => "11110011",
                     30712 => "10100101",
                     30713 => "11110001",
                     30714 => "11010000",
                     30715 => "00011111",
                     30716 => "10101101",
                     30717 => "10110001",
                     30718 => "00000111",
                     30719 => "00101001",
                     30720 => "10010001",
                     30721 => "11010000",
                     30722 => "00001110",
                     30723 => "10101100",
                     30724 => "10110111",
                     30725 => "00000111",
                     30726 => "11110000",
                     30727 => "00000011",
                     30728 => "11001110",
                     30729 => "10110111",
                     30730 => "00000111",
                     30731 => "00100000",
                     30732 => "11110101",
                     30733 => "11111000",
                     30734 => "10001101",
                     30735 => "00000000",
                     30736 => "01000000",
                     30737 => "10101101",
                     30738 => "11001010",
                     30739 => "00000111",
                     30740 => "11010000",
                     30741 => "00000010",
                     30742 => "10101001",
                     30743 => "01111111",
                     30744 => "10001101",
                     30745 => "00000001",
                     30746 => "01000000",
                     30747 => "10100101",
                     30748 => "11111001",
                     30749 => "11001110",
                     30750 => "10111001",
                     30751 => "00000111",
                     30752 => "11010000",
                     30753 => "01001100",
                     30754 => "10100100",
                     30755 => "11111001",
                     30756 => "11100110",
                     30757 => "11111001",
                     30758 => "10110001",
                     30759 => "11110101",
                     30760 => "11110000",
                     30761 => "01000001",
                     30762 => "00010000",
                     30763 => "00010011",
                     30764 => "00100000",
                     30765 => "11001100",
                     30766 => "11111000",
                     30767 => "10001101",
                     30768 => "10111000",
                     30769 => "00000111",
                     30770 => "10101001",
                     30771 => "00011111",
                     30772 => "10001101",
                     30773 => "00001000",
                     30774 => "01000000",
                     30775 => "10100100",
                     30776 => "11111001",
                     30777 => "11100110",
                     30778 => "11111001",
                     30779 => "10110001",
                     30780 => "11110101",
                     30781 => "11110000",
                     30782 => "00101100",
                     30783 => "00100000",
                     30784 => "10101110",
                     30785 => "11110011",
                     30786 => "10101110",
                     30787 => "10111000",
                     30788 => "00000111",
                     30789 => "10001110",
                     30790 => "10111001",
                     30791 => "00000111",
                     30792 => "10101101",
                     30793 => "10110001",
                     30794 => "00000111",
                     30795 => "00101001",
                     30796 => "01101110",
                     30797 => "11010000",
                     30798 => "00000110",
                     30799 => "10100101",
                     30800 => "11110100",
                     30801 => "00101001",
                     30802 => "00001010",
                     30803 => "11110000",
                     30804 => "00011001",
                     30805 => "10001010",
                     30806 => "11001001",
                     30807 => "00010010",
                     30808 => "10110000",
                     30809 => "00001111",
                     30810 => "10101101",
                     30811 => "10110001",
                     30812 => "00000111",
                     30813 => "00101001",
                     30814 => "00001000",
                     30815 => "11110000",
                     30816 => "00000100",
                     30817 => "10101001",
                     30818 => "00001111",
                     30819 => "11010000",
                     30820 => "00000110",
                     30821 => "10101001",
                     30822 => "00011111",
                     30823 => "11010000",
                     30824 => "00000010",
                     30825 => "10101001",
                     30826 => "11111111",
                     30827 => "10001101",
                     30828 => "00001000",
                     30829 => "01000000",
                     30830 => "10100101",
                     30831 => "11110100",
                     30832 => "00101001",
                     30833 => "11110011",
                     30834 => "11110000",
                     30835 => "01010001",
                     30836 => "11001110",
                     30837 => "10111010",
                     30838 => "00000111",
                     30839 => "11010000",
                     30840 => "01001100",
                     30841 => "10101100",
                     30842 => "10110000",
                     30843 => "00000111",
                     30844 => "11101110",
                     30845 => "10110000",
                     30846 => "00000111",
                     30847 => "10110001",
                     30848 => "11110101",
                     30849 => "11010000",
                     30850 => "00001000",
                     30851 => "10101101",
                     30852 => "11000001",
                     30853 => "00000111",
                     30854 => "10001101",
                     30855 => "10110000",
                     30856 => "00000111",
                     30857 => "11010000",
                     30858 => "11101110",
                     30859 => "00100000",
                     30860 => "11000110",
                     30861 => "11111000",
                     30862 => "10001101",
                     30863 => "10111010",
                     30864 => "00000111",
                     30865 => "10001010",
                     30866 => "00101001",
                     30867 => "00111110",
                     30868 => "11110000",
                     30869 => "00100100",
                     30870 => "11001001",
                     30871 => "00110000",
                     30872 => "11110000",
                     30873 => "00011000",
                     30874 => "11001001",
                     30875 => "00100000",
                     30876 => "11110000",
                     30877 => "00001100",
                     30878 => "00101001",
                     30879 => "00010000",
                     30880 => "11110000",
                     30881 => "00011000",
                     30882 => "10101001",
                     30883 => "00011100",
                     30884 => "10100010",
                     30885 => "00000011",
                     30886 => "10100000",
                     30887 => "00011000",
                     30888 => "11010000",
                     30889 => "00010010",
                     30890 => "10101001",
                     30891 => "00011100",
                     30892 => "10100010",
                     30893 => "00001100",
                     30894 => "10100000",
                     30895 => "00011000",
                     30896 => "11010000",
                     30897 => "00001010",
                     30898 => "10101001",
                     30899 => "00011100",
                     30900 => "10100010",
                     30901 => "00000011",
                     30902 => "10100000",
                     30903 => "01011000",
                     30904 => "11010000",
                     30905 => "00000010",
                     30906 => "10101001",
                     30907 => "00010000",
                     30908 => "10001101",
                     30909 => "00001100",
                     30910 => "01000000",
                     30911 => "10001110",
                     30912 => "00001110",
                     30913 => "01000000",
                     30914 => "10001100",
                     30915 => "00001111",
                     30916 => "01000000",
                     30917 => "01100000",
                     30918 => "10101010",
                     30919 => "01101010",
                     30920 => "10001010",
                     30921 => "00101010",
                     30922 => "00101010",
                     30923 => "00101010",
                     30924 => "00101001",
                     30925 => "00000111",
                     30926 => "00011000",
                     30927 => "01100101",
                     30928 => "11110000",
                     30929 => "01101101",
                     30930 => "11000100",
                     30931 => "00000111",
                     30932 => "10101000",
                     30933 => "10111001",
                     30934 => "01100110",
                     30935 => "11111111",
                     30936 => "01100000",
                     30937 => "10101101",
                     30938 => "10110001",
                     30939 => "00000111",
                     30940 => "00101001",
                     30941 => "00001000",
                     30942 => "11110000",
                     30943 => "00000100",
                     30944 => "10101001",
                     30945 => "00000100",
                     30946 => "11010000",
                     30947 => "00001100",
                     30948 => "10100101",
                     30949 => "11110100",
                     30950 => "00101001",
                     30951 => "01111101",
                     30952 => "11110000",
                     30953 => "00000100",
                     30954 => "10101001",
                     30955 => "00001000",
                     30956 => "11010000",
                     30957 => "00000010",
                     30958 => "10101001",
                     30959 => "00101000",
                     30960 => "10100010",
                     30961 => "10000010",
                     30962 => "10100000",
                     30963 => "01111111",
                     30964 => "01100000",
                     30965 => "10101101",
                     30966 => "10110001",
                     30967 => "00000111",
                     30968 => "00101001",
                     30969 => "00001000",
                     30970 => "11110000",
                     30971 => "00000100",
                     30972 => "10111001",
                     30973 => "10010110",
                     30974 => "11111111",
                     30975 => "01100000",
                     30976 => "10100101",
                     30977 => "11110100",
                     30978 => "00101001",
                     30979 => "01111101",
                     30980 => "11110000",
                     30981 => "00000100",
                     30982 => "10111001",
                     30983 => "10011010",
                     30984 => "11111111",
                     30985 => "01100000",
                     30986 => "10111001",
                     30987 => "10100010",
                     30988 => "11111111",
                     30989 => "01100000",
                     30990 => "10100101",
                     30991 => "01011001",
                     30992 => "01010100",
                     30993 => "01100100",
                     30994 => "01011001",
                     30995 => "00111100",
                     30996 => "00110001",
                     30997 => "01001011",
                     30998 => "01101001",
                     30999 => "01011110",
                     31000 => "01000110",
                     31001 => "01001111",
                     31002 => "00110110",
                     31003 => "10001101",
                     31004 => "00110110",
                     31005 => "01001011",
                     31006 => "10001101",
                     31007 => "01101001",
                     31008 => "01101001",
                     31009 => "01101111",
                     31010 => "01110101",
                     31011 => "01101111",
                     31012 => "01111011",
                     31013 => "01101111",
                     31014 => "01110101",
                     31015 => "01101111",
                     31016 => "01111011",
                     31017 => "10000001",
                     31018 => "10000111",
                     31019 => "10000001",
                     31020 => "10001101",
                     31021 => "01101001",
                     31022 => "01101001",
                     31023 => "10010011",
                     31024 => "10011001",
                     31025 => "10010011",
                     31026 => "10011111",
                     31027 => "10010011",
                     31028 => "10011001",
                     31029 => "10010011",
                     31030 => "10011111",
                     31031 => "10000001",
                     31032 => "10000111",
                     31033 => "10000001",
                     31034 => "10001101",
                     31035 => "10010011",
                     31036 => "10011001",
                     31037 => "10010011",
                     31038 => "10011111",
                     31039 => "00001000",
                     31040 => "01110011",
                     31041 => "11111100",
                     31042 => "00100111",
                     31043 => "00011000",
                     31044 => "00100000",
                     31045 => "10111001",
                     31046 => "11111001",
                     31047 => "00101110",
                     31048 => "00011010",
                     31049 => "01000000",
                     31050 => "00100000",
                     31051 => "10110001",
                     31052 => "11111100",
                     31053 => "00111101",
                     31054 => "00100001",
                     31055 => "00100000",
                     31056 => "11000101",
                     31057 => "11111100",
                     31058 => "00111111",
                     31059 => "00011101",
                     31060 => "00011000",
                     31061 => "00010010",
                     31062 => "11111101",
                     31063 => "00000000",
                     31064 => "00000000",
                     31065 => "00001000",
                     31066 => "00011101",
                     31067 => "11111010",
                     31068 => "00000000",
                     31069 => "00000000",
                     31070 => "10100101",
                     31071 => "11111011",
                     31072 => "10010011",
                     31073 => "01100010",
                     31074 => "00010000",
                     31075 => "11001001",
                     31076 => "11111110",
                     31077 => "00100100",
                     31078 => "00010100",
                     31079 => "00011000",
                     31080 => "01000110",
                     31081 => "11111100",
                     31082 => "00011110",
                     31083 => "00010100",
                     31084 => "00001000",
                     31085 => "01010011",
                     31086 => "11111101",
                     31087 => "10100000",
                     31088 => "01110000",
                     31089 => "01101000",
                     31090 => "00001000",
                     31091 => "01010010",
                     31092 => "11111110",
                     31093 => "01001100",
                     31094 => "00100100",
                     31095 => "00011000",
                     31096 => "00000010",
                     31097 => "11111010",
                     31098 => "00101101",
                     31099 => "00011100",
                     31100 => "10111000",
                     31101 => "00011000",
                     31102 => "01001010",
                     31103 => "11111010",
                     31104 => "00100000",
                     31105 => "00010010",
                     31106 => "01110000",
                     31107 => "00011000",
                     31108 => "01110110",
                     31109 => "11111010",
                     31110 => "00011011",
                     31111 => "00010000",
                     31112 => "01000100",
                     31113 => "00011000",
                     31114 => "10011110",
                     31115 => "11111010",
                     31116 => "00010001",
                     31117 => "00001010",
                     31118 => "00011100",
                     31119 => "00011000",
                     31120 => "11000011",
                     31121 => "11111010",
                     31122 => "00101101",
                     31123 => "00010000",
                     31124 => "01011000",
                     31125 => "00011000",
                     31126 => "11011100",
                     31127 => "11111010",
                     31128 => "00010100",
                     31129 => "00001101",
                     31130 => "00111111",
                     31131 => "00011000",
                     31132 => "11111010",
                     31133 => "11111010",
                     31134 => "00010101",
                     31135 => "00001101",
                     31136 => "00100001",
                     31137 => "00011000",
                     31138 => "00100110",
                     31139 => "11111011",
                     31140 => "00011000",
                     31141 => "00010000",
                     31142 => "01111010",
                     31143 => "00011000",
                     31144 => "01001100",
                     31145 => "11111011",
                     31146 => "00011001",
                     31147 => "00001111",
                     31148 => "01010100",
                     31149 => "00011000",
                     31150 => "01110101",
                     31151 => "11111011",
                     31152 => "00011110",
                     31153 => "00010010",
                     31154 => "00101011",
                     31155 => "00011000",
                     31156 => "01110011",
                     31157 => "11111011",
                     31158 => "00011110",
                     31159 => "00001111",
                     31160 => "00101101",
                     31161 => "10000100",
                     31162 => "00101100",
                     31163 => "00101100",
                     31164 => "00101100",
                     31165 => "10000010",
                     31166 => "00000100",
                     31167 => "00101100",
                     31168 => "00000100",
                     31169 => "10000101",
                     31170 => "00101100",
                     31171 => "10000100",
                     31172 => "00101100",
                     31173 => "00101100",
                     31174 => "00101010",
                     31175 => "00101010",
                     31176 => "00101010",
                     31177 => "10000010",
                     31178 => "00000100",
                     31179 => "00101010",
                     31180 => "00000100",
                     31181 => "10000101",
                     31182 => "00101010",
                     31183 => "10000100",
                     31184 => "00101010",
                     31185 => "00101010",
                     31186 => "00000000",
                     31187 => "00011111",
                     31188 => "00011111",
                     31189 => "00011111",
                     31190 => "10011000",
                     31191 => "00011111",
                     31192 => "00011111",
                     31193 => "10011000",
                     31194 => "10011110",
                     31195 => "10011000",
                     31196 => "00011111",
                     31197 => "00011101",
                     31198 => "00011101",
                     31199 => "00011101",
                     31200 => "10010100",
                     31201 => "00011101",
                     31202 => "00011101",
                     31203 => "10010100",
                     31204 => "10011100",
                     31205 => "10010100",
                     31206 => "00011101",
                     31207 => "10000110",
                     31208 => "00011000",
                     31209 => "10000101",
                     31210 => "00100110",
                     31211 => "00110000",
                     31212 => "10000100",
                     31213 => "00000100",
                     31214 => "00100110",
                     31215 => "00110000",
                     31216 => "10000110",
                     31217 => "00010100",
                     31218 => "10000101",
                     31219 => "00100010",
                     31220 => "00101100",
                     31221 => "10000100",
                     31222 => "00000100",
                     31223 => "00100010",
                     31224 => "00101100",
                     31225 => "00100001",
                     31226 => "11010000",
                     31227 => "11000100",
                     31228 => "11010000",
                     31229 => "00110001",
                     31230 => "11010000",
                     31231 => "11000100",
                     31232 => "11010000",
                     31233 => "00000000",
                     31234 => "10000101",
                     31235 => "00101100",
                     31236 => "00100010",
                     31237 => "00011100",
                     31238 => "10000100",
                     31239 => "00100110",
                     31240 => "00101010",
                     31241 => "10000010",
                     31242 => "00101000",
                     31243 => "00100110",
                     31244 => "00000100",
                     31245 => "10000111",
                     31246 => "00100010",
                     31247 => "00110100",
                     31248 => "00111010",
                     31249 => "10000010",
                     31250 => "01000000",
                     31251 => "00000100",
                     31252 => "00110110",
                     31253 => "10000100",
                     31254 => "00111010",
                     31255 => "00110100",
                     31256 => "10000010",
                     31257 => "00101100",
                     31258 => "00110000",
                     31259 => "10000101",
                     31260 => "00101010",
                     31261 => "00000000",
                     31262 => "01011101",
                     31263 => "01010101",
                     31264 => "01001101",
                     31265 => "00010101",
                     31266 => "00011001",
                     31267 => "10010110",
                     31268 => "00010101",
                     31269 => "11010101",
                     31270 => "11100011",
                     31271 => "11101011",
                     31272 => "00101101",
                     31273 => "10100110",
                     31274 => "00101011",
                     31275 => "00100111",
                     31276 => "10011100",
                     31277 => "10011110",
                     31278 => "01011001",
                     31279 => "10000101",
                     31280 => "00100010",
                     31281 => "00011100",
                     31282 => "00010100",
                     31283 => "10000100",
                     31284 => "00011110",
                     31285 => "00100010",
                     31286 => "10000010",
                     31287 => "00100000",
                     31288 => "00011110",
                     31289 => "00000100",
                     31290 => "10000111",
                     31291 => "00011100",
                     31292 => "00101100",
                     31293 => "00110100",
                     31294 => "10000010",
                     31295 => "00110110",
                     31296 => "00000100",
                     31297 => "00110000",
                     31298 => "00110100",
                     31299 => "00000100",
                     31300 => "00101100",
                     31301 => "00000100",
                     31302 => "00100110",
                     31303 => "00101010",
                     31304 => "10000101",
                     31305 => "00100010",
                     31306 => "10000100",
                     31307 => "00000100",
                     31308 => "10000010",
                     31309 => "00111010",
                     31310 => "00111000",
                     31311 => "00110110",
                     31312 => "00110010",
                     31313 => "00000100",
                     31314 => "00110100",
                     31315 => "00000100",
                     31316 => "00100100",
                     31317 => "00100110",
                     31318 => "00101100",
                     31319 => "00000100",
                     31320 => "00100110",
                     31321 => "00101100",
                     31322 => "00110000",
                     31323 => "00000000",
                     31324 => "00000101",
                     31325 => "10110100",
                     31326 => "10110010",
                     31327 => "10110000",
                     31328 => "00101011",
                     31329 => "10101100",
                     31330 => "10000100",
                     31331 => "10011100",
                     31332 => "10011110",
                     31333 => "10100010",
                     31334 => "10000100",
                     31335 => "10010100",
                     31336 => "10011100",
                     31337 => "10011110",
                     31338 => "10000101",
                     31339 => "00010100",
                     31340 => "00100010",
                     31341 => "10000100",
                     31342 => "00101100",
                     31343 => "10000101",
                     31344 => "00011110",
                     31345 => "10000010",
                     31346 => "00101100",
                     31347 => "10000100",
                     31348 => "00101100",
                     31349 => "00011110",
                     31350 => "10000100",
                     31351 => "00000100",
                     31352 => "10000010",
                     31353 => "00111010",
                     31354 => "00111000",
                     31355 => "00110110",
                     31356 => "00110010",
                     31357 => "00000100",
                     31358 => "00110100",
                     31359 => "00000100",
                     31360 => "01100100",
                     31361 => "00000100",
                     31362 => "01100100",
                     31363 => "10000110",
                     31364 => "01100100",
                     31365 => "00000000",
                     31366 => "00000101",
                     31367 => "10110100",
                     31368 => "10110010",
                     31369 => "10110000",
                     31370 => "00101011",
                     31371 => "10101100",
                     31372 => "10000100",
                     31373 => "00110111",
                     31374 => "10110110",
                     31375 => "10110110",
                     31376 => "01000101",
                     31377 => "10000101",
                     31378 => "00010100",
                     31379 => "00011100",
                     31380 => "10000010",
                     31381 => "00100010",
                     31382 => "10000100",
                     31383 => "00101100",
                     31384 => "01001110",
                     31385 => "10000010",
                     31386 => "01001110",
                     31387 => "10000100",
                     31388 => "01001110",
                     31389 => "00100010",
                     31390 => "10000100",
                     31391 => "00000100",
                     31392 => "10000101",
                     31393 => "00110010",
                     31394 => "10000101",
                     31395 => "00110000",
                     31396 => "10000110",
                     31397 => "00101100",
                     31398 => "00000100",
                     31399 => "00000000",
                     31400 => "00000101",
                     31401 => "10100100",
                     31402 => "00000101",
                     31403 => "10011110",
                     31404 => "00000101",
                     31405 => "10011101",
                     31406 => "10000101",
                     31407 => "10000100",
                     31408 => "00010100",
                     31409 => "10000101",
                     31410 => "00100100",
                     31411 => "00101000",
                     31412 => "00101100",
                     31413 => "10000010",
                     31414 => "00100010",
                     31415 => "10000100",
                     31416 => "00100010",
                     31417 => "00010100",
                     31418 => "00100001",
                     31419 => "11010000",
                     31420 => "11000100",
                     31421 => "11010000",
                     31422 => "00110001",
                     31423 => "11010000",
                     31424 => "11000100",
                     31425 => "11010000",
                     31426 => "00000000",
                     31427 => "10000010",
                     31428 => "00101100",
                     31429 => "10000100",
                     31430 => "00101100",
                     31431 => "00101100",
                     31432 => "10000010",
                     31433 => "00101100",
                     31434 => "00110000",
                     31435 => "00000100",
                     31436 => "00110100",
                     31437 => "00101100",
                     31438 => "00000100",
                     31439 => "00100110",
                     31440 => "10000110",
                     31441 => "00100010",
                     31442 => "00000000",
                     31443 => "10100100",
                     31444 => "00100101",
                     31445 => "00100101",
                     31446 => "10100100",
                     31447 => "00101001",
                     31448 => "10100010",
                     31449 => "00011101",
                     31450 => "10011100",
                     31451 => "10010101",
                     31452 => "10000010",
                     31453 => "00101100",
                     31454 => "00101100",
                     31455 => "00000100",
                     31456 => "00101100",
                     31457 => "00000100",
                     31458 => "00101100",
                     31459 => "00110000",
                     31460 => "10000101",
                     31461 => "00110100",
                     31462 => "00000100",
                     31463 => "00000100",
                     31464 => "00000000",
                     31465 => "10100100",
                     31466 => "00100101",
                     31467 => "00100101",
                     31468 => "10100100",
                     31469 => "10101000",
                     31470 => "01100011",
                     31471 => "00000100",
                     31472 => "10000101",
                     31473 => "00001110",
                     31474 => "00011010",
                     31475 => "10000100",
                     31476 => "00100100",
                     31477 => "10000101",
                     31478 => "00100010",
                     31479 => "00010100",
                     31480 => "10000100",
                     31481 => "00001100",
                     31482 => "10000010",
                     31483 => "00110100",
                     31484 => "10000100",
                     31485 => "00110100",
                     31486 => "00110100",
                     31487 => "10000010",
                     31488 => "00101100",
                     31489 => "10000100",
                     31490 => "00110100",
                     31491 => "10000110",
                     31492 => "00111010",
                     31493 => "00000100",
                     31494 => "00000000",
                     31495 => "10100000",
                     31496 => "00100001",
                     31497 => "00100001",
                     31498 => "10100000",
                     31499 => "00100001",
                     31500 => "00101011",
                     31501 => "00000101",
                     31502 => "10100011",
                     31503 => "10000010",
                     31504 => "00011000",
                     31505 => "10000100",
                     31506 => "00011000",
                     31507 => "00011000",
                     31508 => "10000010",
                     31509 => "00011000",
                     31510 => "00011000",
                     31511 => "00000100",
                     31512 => "10000110",
                     31513 => "00111010",
                     31514 => "00100010",
                     31515 => "00110001",
                     31516 => "10010000",
                     31517 => "00110001",
                     31518 => "10010000",
                     31519 => "00110001",
                     31520 => "01110001",
                     31521 => "00110001",
                     31522 => "10010000",
                     31523 => "10010000",
                     31524 => "10010000",
                     31525 => "00000000",
                     31526 => "10000010",
                     31527 => "00110100",
                     31528 => "10000100",
                     31529 => "00101100",
                     31530 => "10000101",
                     31531 => "00100010",
                     31532 => "10000100",
                     31533 => "00100100",
                     31534 => "10000010",
                     31535 => "00100110",
                     31536 => "00110110",
                     31537 => "00000100",
                     31538 => "00110110",
                     31539 => "10000110",
                     31540 => "00100110",
                     31541 => "00000000",
                     31542 => "10101100",
                     31543 => "00100111",
                     31544 => "01011101",
                     31545 => "00011101",
                     31546 => "10011110",
                     31547 => "00101101",
                     31548 => "10101100",
                     31549 => "10011111",
                     31550 => "10000101",
                     31551 => "00010100",
                     31552 => "10000010",
                     31553 => "00100000",
                     31554 => "10000100",
                     31555 => "00100010",
                     31556 => "00101100",
                     31557 => "00011110",
                     31558 => "00011110",
                     31559 => "10000010",
                     31560 => "00101100",
                     31561 => "00101100",
                     31562 => "00011110",
                     31563 => "00000100",
                     31564 => "10000111",
                     31565 => "00101010",
                     31566 => "01000000",
                     31567 => "01000000",
                     31568 => "01000000",
                     31569 => "00111010",
                     31570 => "00110110",
                     31571 => "10000010",
                     31572 => "00110100",
                     31573 => "00101100",
                     31574 => "00000100",
                     31575 => "00100110",
                     31576 => "10000110",
                     31577 => "00100010",
                     31578 => "00000000",
                     31579 => "11100011",
                     31580 => "11110111",
                     31581 => "11110111",
                     31582 => "11110111",
                     31583 => "11110101",
                     31584 => "11110001",
                     31585 => "10101100",
                     31586 => "00100111",
                     31587 => "10011110",
                     31588 => "10011101",
                     31589 => "10000101",
                     31590 => "00011000",
                     31591 => "10000010",
                     31592 => "00011110",
                     31593 => "10000100",
                     31594 => "00100010",
                     31595 => "00101010",
                     31596 => "00100010",
                     31597 => "00100010",
                     31598 => "10000010",
                     31599 => "00101100",
                     31600 => "00101100",
                     31601 => "00100010",
                     31602 => "00000100",
                     31603 => "10000110",
                     31604 => "00000100",
                     31605 => "10000010",
                     31606 => "00101010",
                     31607 => "00110110",
                     31608 => "00000100",
                     31609 => "00110110",
                     31610 => "10000111",
                     31611 => "00110110",
                     31612 => "00110100",
                     31613 => "00110000",
                     31614 => "10000110",
                     31615 => "00101100",
                     31616 => "00000100",
                     31617 => "00000000",
                     31618 => "00000000",
                     31619 => "01101000",
                     31620 => "01101010",
                     31621 => "01101100",
                     31622 => "01000101",
                     31623 => "10100010",
                     31624 => "00110001",
                     31625 => "10110000",
                     31626 => "11110001",
                     31627 => "11101101",
                     31628 => "11101011",
                     31629 => "10100010",
                     31630 => "00011101",
                     31631 => "10011100",
                     31632 => "10010101",
                     31633 => "10000110",
                     31634 => "00000100",
                     31635 => "10000101",
                     31636 => "00100010",
                     31637 => "10000010",
                     31638 => "00100010",
                     31639 => "10000111",
                     31640 => "00100010",
                     31641 => "00100110",
                     31642 => "00101010",
                     31643 => "10000100",
                     31644 => "00101100",
                     31645 => "00100010",
                     31646 => "10000110",
                     31647 => "00010100",
                     31648 => "01010001",
                     31649 => "10010000",
                     31650 => "00110001",
                     31651 => "00010001",
                     31652 => "00000000",
                     31653 => "10000000",
                     31654 => "00100010",
                     31655 => "00101000",
                     31656 => "00100010",
                     31657 => "00100110",
                     31658 => "00100010",
                     31659 => "00100100",
                     31660 => "00100010",
                     31661 => "00100110",
                     31662 => "00100010",
                     31663 => "00101000",
                     31664 => "00100010",
                     31665 => "00101010",
                     31666 => "00100010",
                     31667 => "00101000",
                     31668 => "00100010",
                     31669 => "00100110",
                     31670 => "00100010",
                     31671 => "00101000",
                     31672 => "00100010",
                     31673 => "00100110",
                     31674 => "00100010",
                     31675 => "00100100",
                     31676 => "00100010",
                     31677 => "00100110",
                     31678 => "00100010",
                     31679 => "00101000",
                     31680 => "00100010",
                     31681 => "00101010",
                     31682 => "00100010",
                     31683 => "00101000",
                     31684 => "00100010",
                     31685 => "00100110",
                     31686 => "00100000",
                     31687 => "00100110",
                     31688 => "00100000",
                     31689 => "00100100",
                     31690 => "00100000",
                     31691 => "00100110",
                     31692 => "00100000",
                     31693 => "00101000",
                     31694 => "00100000",
                     31695 => "00100110",
                     31696 => "00100000",
                     31697 => "00101000",
                     31698 => "00100000",
                     31699 => "00100110",
                     31700 => "00100000",
                     31701 => "00100100",
                     31702 => "00100000",
                     31703 => "00100110",
                     31704 => "00100000",
                     31705 => "00100100",
                     31706 => "00100000",
                     31707 => "00100110",
                     31708 => "00100000",
                     31709 => "00101000",
                     31710 => "00100000",
                     31711 => "00100110",
                     31712 => "00100000",
                     31713 => "00101000",
                     31714 => "00100000",
                     31715 => "00100110",
                     31716 => "00100000",
                     31717 => "00100100",
                     31718 => "00101000",
                     31719 => "00110000",
                     31720 => "00101000",
                     31721 => "00110010",
                     31722 => "00101000",
                     31723 => "00110000",
                     31724 => "00101000",
                     31725 => "00101110",
                     31726 => "00101000",
                     31727 => "00110000",
                     31728 => "00101000",
                     31729 => "00101110",
                     31730 => "00101000",
                     31731 => "00101100",
                     31732 => "00101000",
                     31733 => "00101110",
                     31734 => "00101000",
                     31735 => "00110000",
                     31736 => "00101000",
                     31737 => "00110010",
                     31738 => "00101000",
                     31739 => "00110000",
                     31740 => "00101000",
                     31741 => "00101110",
                     31742 => "00101000",
                     31743 => "00110000",
                     31744 => "00101000",
                     31745 => "00101110",
                     31746 => "00101000",
                     31747 => "00101100",
                     31748 => "00101000",
                     31749 => "00101110",
                     31750 => "00000000",
                     31751 => "00000100",
                     31752 => "01110000",
                     31753 => "01101110",
                     31754 => "01101100",
                     31755 => "01101110",
                     31756 => "01110000",
                     31757 => "01110010",
                     31758 => "01110000",
                     31759 => "01101110",
                     31760 => "01110000",
                     31761 => "01101110",
                     31762 => "01101100",
                     31763 => "01101110",
                     31764 => "01110000",
                     31765 => "01110010",
                     31766 => "01110000",
                     31767 => "01101110",
                     31768 => "01101110",
                     31769 => "01101100",
                     31770 => "01101110",
                     31771 => "01110000",
                     31772 => "01101110",
                     31773 => "01110000",
                     31774 => "01101110",
                     31775 => "01101100",
                     31776 => "01101110",
                     31777 => "01101100",
                     31778 => "01101110",
                     31779 => "01110000",
                     31780 => "01101110",
                     31781 => "01110000",
                     31782 => "01101110",
                     31783 => "01101100",
                     31784 => "01110110",
                     31785 => "01111000",
                     31786 => "01110110",
                     31787 => "01110100",
                     31788 => "01110110",
                     31789 => "01110100",
                     31790 => "01110010",
                     31791 => "01110100",
                     31792 => "01110110",
                     31793 => "01111000",
                     31794 => "01110110",
                     31795 => "01110100",
                     31796 => "01110110",
                     31797 => "01110100",
                     31798 => "01110010",
                     31799 => "01110100",
                     31800 => "10000100",
                     31801 => "00011010",
                     31802 => "10000011",
                     31803 => "00011000",
                     31804 => "00100000",
                     31805 => "10000100",
                     31806 => "00011110",
                     31807 => "10000011",
                     31808 => "00011100",
                     31809 => "00101000",
                     31810 => "00100110",
                     31811 => "00011100",
                     31812 => "00011010",
                     31813 => "00011100",
                     31814 => "10000010",
                     31815 => "00101100",
                     31816 => "00000100",
                     31817 => "00000100",
                     31818 => "00100010",
                     31819 => "00000100",
                     31820 => "00000100",
                     31821 => "10000100",
                     31822 => "00011100",
                     31823 => "10000111",
                     31824 => "00100110",
                     31825 => "00101010",
                     31826 => "00100110",
                     31827 => "10000100",
                     31828 => "00100100",
                     31829 => "00101000",
                     31830 => "00100100",
                     31831 => "10000000",
                     31832 => "00100010",
                     31833 => "00000000",
                     31834 => "10011100",
                     31835 => "00000101",
                     31836 => "10010100",
                     31837 => "00000101",
                     31838 => "00001101",
                     31839 => "10011111",
                     31840 => "00011110",
                     31841 => "10011100",
                     31842 => "10011000",
                     31843 => "10011101",
                     31844 => "10000010",
                     31845 => "00100010",
                     31846 => "00000100",
                     31847 => "00000100",
                     31848 => "00011100",
                     31849 => "00000100",
                     31850 => "00000100",
                     31851 => "10000100",
                     31852 => "00010100",
                     31853 => "10000110",
                     31854 => "00011110",
                     31855 => "10000000",
                     31856 => "00010110",
                     31857 => "10000000",
                     31858 => "00010100",
                     31859 => "10000001",
                     31860 => "00011100",
                     31861 => "00110000",
                     31862 => "00000100",
                     31863 => "00110000",
                     31864 => "00110000",
                     31865 => "00000100",
                     31866 => "00011110",
                     31867 => "00110010",
                     31868 => "00000100",
                     31869 => "00110010",
                     31870 => "00110010",
                     31871 => "00000100",
                     31872 => "00100000",
                     31873 => "00110100",
                     31874 => "00000100",
                     31875 => "00110100",
                     31876 => "00110100",
                     31877 => "00000100",
                     31878 => "00110110",
                     31879 => "00000100",
                     31880 => "10000100",
                     31881 => "00110110",
                     31882 => "00000000",
                     31883 => "01000110",
                     31884 => "10100100",
                     31885 => "01100100",
                     31886 => "10100100",
                     31887 => "01001000",
                     31888 => "10100110",
                     31889 => "01100110",
                     31890 => "10100110",
                     31891 => "01001010",
                     31892 => "10101000",
                     31893 => "01101000",
                     31894 => "10101000",
                     31895 => "01101010",
                     31896 => "01000100",
                     31897 => "00101011",
                     31898 => "10000001",
                     31899 => "00101010",
                     31900 => "01000010",
                     31901 => "00000100",
                     31902 => "01000010",
                     31903 => "01000010",
                     31904 => "00000100",
                     31905 => "00101100",
                     31906 => "01100100",
                     31907 => "00000100",
                     31908 => "01100100",
                     31909 => "01100100",
                     31910 => "00000100",
                     31911 => "00101110",
                     31912 => "01000110",
                     31913 => "00000100",
                     31914 => "01000110",
                     31915 => "01000110",
                     31916 => "00000100",
                     31917 => "00100010",
                     31918 => "00000100",
                     31919 => "10000100",
                     31920 => "00100010",
                     31921 => "10000111",
                     31922 => "00000100",
                     31923 => "00000110",
                     31924 => "00001100",
                     31925 => "00010100",
                     31926 => "00011100",
                     31927 => "00100010",
                     31928 => "10000110",
                     31929 => "00101100",
                     31930 => "00100010",
                     31931 => "10000111",
                     31932 => "00000100",
                     31933 => "01100000",
                     31934 => "00001110",
                     31935 => "00010100",
                     31936 => "00011010",
                     31937 => "00100100",
                     31938 => "10000110",
                     31939 => "00101100",
                     31940 => "00100100",
                     31941 => "10000111",
                     31942 => "00000100",
                     31943 => "00001000",
                     31944 => "00010000",
                     31945 => "00011000",
                     31946 => "00011110",
                     31947 => "00101000",
                     31948 => "10000110",
                     31949 => "00110000",
                     31950 => "00110000",
                     31951 => "10000000",
                     31952 => "01100100",
                     31953 => "00000000",
                     31954 => "11001101",
                     31955 => "11010101",
                     31956 => "11011101",
                     31957 => "11100011",
                     31958 => "11101101",
                     31959 => "11110101",
                     31960 => "10111011",
                     31961 => "10110101",
                     31962 => "11001111",
                     31963 => "11010101",
                     31964 => "11011011",
                     31965 => "11100101",
                     31966 => "11101101",
                     31967 => "11110011",
                     31968 => "10111101",
                     31969 => "10110011",
                     31970 => "11010001",
                     31971 => "11011001",
                     31972 => "11011111",
                     31973 => "11101001",
                     31974 => "11110001",
                     31975 => "11110111",
                     31976 => "10111111",
                     31977 => "11111111",
                     31978 => "11111111",
                     31979 => "11111111",
                     31980 => "00110100",
                     31981 => "00000000",
                     31982 => "10000110",
                     31983 => "00000100",
                     31984 => "10000111",
                     31985 => "00010100",
                     31986 => "00011100",
                     31987 => "00100010",
                     31988 => "10000110",
                     31989 => "00110100",
                     31990 => "10000100",
                     31991 => "00101100",
                     31992 => "00000100",
                     31993 => "00000100",
                     31994 => "00000100",
                     31995 => "10000111",
                     31996 => "00010100",
                     31997 => "00011010",
                     31998 => "00100100",
                     31999 => "10000110",
                     32000 => "00110010",
                     32001 => "10000100",
                     32002 => "00101100",
                     32003 => "00000100",
                     32004 => "10000110",
                     32005 => "00000100",
                     32006 => "10000111",
                     32007 => "00011000",
                     32008 => "00011110",
                     32009 => "00101000",
                     32010 => "10000110",
                     32011 => "00110110",
                     32012 => "10000111",
                     32013 => "00110000",
                     32014 => "00110000",
                     32015 => "00110000",
                     32016 => "10000000",
                     32017 => "00101100",
                     32018 => "10000010",
                     32019 => "00010100",
                     32020 => "00101100",
                     32021 => "01100010",
                     32022 => "00100110",
                     32023 => "00010000",
                     32024 => "00101000",
                     32025 => "10000000",
                     32026 => "00000100",
                     32027 => "10000010",
                     32028 => "00010100",
                     32029 => "00101100",
                     32030 => "01100010",
                     32031 => "00100110",
                     32032 => "00010000",
                     32033 => "00101000",
                     32034 => "10000000",
                     32035 => "00000100",
                     32036 => "10000010",
                     32037 => "00001000",
                     32038 => "00011110",
                     32039 => "01011110",
                     32040 => "00011000",
                     32041 => "01100000",
                     32042 => "00011010",
                     32043 => "10000000",
                     32044 => "00000100",
                     32045 => "10000010",
                     32046 => "00001000",
                     32047 => "00011110",
                     32048 => "01011110",
                     32049 => "00011000",
                     32050 => "01100000",
                     32051 => "00011010",
                     32052 => "10000110",
                     32053 => "00000100",
                     32054 => "10000011",
                     32055 => "00011010",
                     32056 => "00011000",
                     32057 => "00010110",
                     32058 => "10000100",
                     32059 => "00010100",
                     32060 => "00011010",
                     32061 => "00011000",
                     32062 => "00001110",
                     32063 => "00001100",
                     32064 => "00010110",
                     32065 => "10000011",
                     32066 => "00010100",
                     32067 => "00100000",
                     32068 => "00011110",
                     32069 => "00011100",
                     32070 => "00101000",
                     32071 => "00100110",
                     32072 => "10000111",
                     32073 => "00100100",
                     32074 => "00011010",
                     32075 => "00010010",
                     32076 => "00010000",
                     32077 => "01100010",
                     32078 => "00001110",
                     32079 => "10000000",
                     32080 => "00000100",
                     32081 => "00000100",
                     32082 => "00000000",
                     32083 => "10000010",
                     32084 => "00011000",
                     32085 => "00011100",
                     32086 => "00100000",
                     32087 => "00100010",
                     32088 => "00100110",
                     32089 => "00101000",
                     32090 => "10000001",
                     32091 => "00101010",
                     32092 => "00101010",
                     32093 => "00101010",
                     32094 => "00000100",
                     32095 => "00101010",
                     32096 => "00000100",
                     32097 => "10000011",
                     32098 => "00101010",
                     32099 => "10000010",
                     32100 => "00100010",
                     32101 => "10000110",
                     32102 => "00110100",
                     32103 => "00110010",
                     32104 => "00110100",
                     32105 => "10000001",
                     32106 => "00000100",
                     32107 => "00100010",
                     32108 => "00100110",
                     32109 => "00101010",
                     32110 => "00101100",
                     32111 => "00110000",
                     32112 => "10000110",
                     32113 => "00110100",
                     32114 => "10000011",
                     32115 => "00110010",
                     32116 => "10000010",
                     32117 => "00110110",
                     32118 => "10000100",
                     32119 => "00110100",
                     32120 => "10000101",
                     32121 => "00000100",
                     32122 => "10000001",
                     32123 => "00100010",
                     32124 => "10000110",
                     32125 => "00110000",
                     32126 => "00101110",
                     32127 => "00110000",
                     32128 => "10000001",
                     32129 => "00000100",
                     32130 => "00100010",
                     32131 => "00100110",
                     32132 => "00101010",
                     32133 => "00101100",
                     32134 => "00101110",
                     32135 => "10000110",
                     32136 => "00110000",
                     32137 => "10000011",
                     32138 => "00100010",
                     32139 => "10000010",
                     32140 => "00110110",
                     32141 => "10000100",
                     32142 => "00110100",
                     32143 => "10000101",
                     32144 => "00000100",
                     32145 => "10000001",
                     32146 => "00100010",
                     32147 => "10000110",
                     32148 => "00111010",
                     32149 => "00111010",
                     32150 => "00111010",
                     32151 => "10000010",
                     32152 => "00111010",
                     32153 => "10000001",
                     32154 => "01000000",
                     32155 => "10000010",
                     32156 => "00000100",
                     32157 => "10000001",
                     32158 => "00111010",
                     32159 => "10000110",
                     32160 => "00110110",
                     32161 => "00110110",
                     32162 => "00110110",
                     32163 => "10000010",
                     32164 => "00110110",
                     32165 => "10000001",
                     32166 => "00111010",
                     32167 => "10000010",
                     32168 => "00000100",
                     32169 => "10000001",
                     32170 => "00110110",
                     32171 => "10000110",
                     32172 => "00110100",
                     32173 => "10000010",
                     32174 => "00100110",
                     32175 => "00101010",
                     32176 => "00110110",
                     32177 => "10000001",
                     32178 => "00110100",
                     32179 => "00110100",
                     32180 => "10000101",
                     32181 => "00110100",
                     32182 => "10000001",
                     32183 => "00101010",
                     32184 => "10000110",
                     32185 => "00101100",
                     32186 => "00000000",
                     32187 => "10000100",
                     32188 => "10010000",
                     32189 => "10110000",
                     32190 => "10000100",
                     32191 => "01010000",
                     32192 => "01010000",
                     32193 => "10110000",
                     32194 => "00000000",
                     32195 => "10011000",
                     32196 => "10010110",
                     32197 => "10010100",
                     32198 => "10010010",
                     32199 => "10010100",
                     32200 => "10010110",
                     32201 => "01011000",
                     32202 => "01011000",
                     32203 => "01011000",
                     32204 => "01000100",
                     32205 => "01011100",
                     32206 => "01000100",
                     32207 => "10011111",
                     32208 => "10100011",
                     32209 => "10100001",
                     32210 => "10100011",
                     32211 => "10000101",
                     32212 => "10100011",
                     32213 => "11100000",
                     32214 => "10100110",
                     32215 => "00100011",
                     32216 => "11000100",
                     32217 => "10011111",
                     32218 => "10011101",
                     32219 => "10011111",
                     32220 => "10000101",
                     32221 => "10011111",
                     32222 => "11010010",
                     32223 => "10100110",
                     32224 => "00100011",
                     32225 => "11000100",
                     32226 => "10110101",
                     32227 => "10110001",
                     32228 => "10101111",
                     32229 => "10000101",
                     32230 => "10110001",
                     32231 => "10101111",
                     32232 => "10101101",
                     32233 => "10000101",
                     32234 => "10010101",
                     32235 => "10011110",
                     32236 => "10100010",
                     32237 => "10101010",
                     32238 => "01101010",
                     32239 => "01101010",
                     32240 => "01101011",
                     32241 => "01011110",
                     32242 => "10011101",
                     32243 => "10000100",
                     32244 => "00000100",
                     32245 => "00000100",
                     32246 => "10000010",
                     32247 => "00100010",
                     32248 => "10000110",
                     32249 => "00100010",
                     32250 => "10000010",
                     32251 => "00010100",
                     32252 => "00100010",
                     32253 => "00101100",
                     32254 => "00010010",
                     32255 => "00100010",
                     32256 => "00101010",
                     32257 => "00010100",
                     32258 => "00100010",
                     32259 => "00101100",
                     32260 => "00011100",
                     32261 => "00100010",
                     32262 => "00101100",
                     32263 => "00010100",
                     32264 => "00100010",
                     32265 => "00101100",
                     32266 => "00010010",
                     32267 => "00100010",
                     32268 => "00101010",
                     32269 => "00010100",
                     32270 => "00100010",
                     32271 => "00101100",
                     32272 => "00011100",
                     32273 => "00100010",
                     32274 => "00101100",
                     32275 => "00011000",
                     32276 => "00100010",
                     32277 => "00101010",
                     32278 => "00010110",
                     32279 => "00100000",
                     32280 => "00101000",
                     32281 => "00011000",
                     32282 => "00100010",
                     32283 => "00101010",
                     32284 => "00010010",
                     32285 => "00100010",
                     32286 => "00101010",
                     32287 => "00011000",
                     32288 => "00100010",
                     32289 => "00101010",
                     32290 => "00010010",
                     32291 => "00100010",
                     32292 => "00101010",
                     32293 => "00010100",
                     32294 => "00100010",
                     32295 => "00101100",
                     32296 => "00001100",
                     32297 => "00100010",
                     32298 => "00101100",
                     32299 => "00010100",
                     32300 => "00100010",
                     32301 => "00110100",
                     32302 => "00010010",
                     32303 => "00100010",
                     32304 => "00110000",
                     32305 => "00010000",
                     32306 => "00100010",
                     32307 => "00101110",
                     32308 => "00010110",
                     32309 => "00100010",
                     32310 => "00110100",
                     32311 => "00011000",
                     32312 => "00100110",
                     32313 => "00110110",
                     32314 => "00010110",
                     32315 => "00100110",
                     32316 => "00110110",
                     32317 => "00010100",
                     32318 => "00100110",
                     32319 => "00110110",
                     32320 => "00010010",
                     32321 => "00100010",
                     32322 => "00110110",
                     32323 => "01011100",
                     32324 => "00100010",
                     32325 => "00110100",
                     32326 => "00001100",
                     32327 => "00100010",
                     32328 => "00100010",
                     32329 => "10000001",
                     32330 => "00011110",
                     32331 => "00011110",
                     32332 => "10000101",
                     32333 => "00011110",
                     32334 => "10000001",
                     32335 => "00010010",
                     32336 => "10000110",
                     32337 => "00010100",
                     32338 => "10000001",
                     32339 => "00101100",
                     32340 => "00100010",
                     32341 => "00011100",
                     32342 => "00101100",
                     32343 => "00100010",
                     32344 => "00011100",
                     32345 => "10000101",
                     32346 => "00101100",
                     32347 => "00000100",
                     32348 => "10000001",
                     32349 => "00101110",
                     32350 => "00100100",
                     32351 => "00011110",
                     32352 => "00101110",
                     32353 => "00100100",
                     32354 => "00011110",
                     32355 => "10000101",
                     32356 => "00101110",
                     32357 => "00000100",
                     32358 => "10000001",
                     32359 => "00110010",
                     32360 => "00101000",
                     32361 => "00100010",
                     32362 => "00110010",
                     32363 => "00101000",
                     32364 => "00100010",
                     32365 => "10000101",
                     32366 => "00110010",
                     32367 => "10000111",
                     32368 => "00110110",
                     32369 => "00110110",
                     32370 => "00110110",
                     32371 => "10000100",
                     32372 => "00111010",
                     32373 => "00000000",
                     32374 => "01011100",
                     32375 => "01010100",
                     32376 => "01001100",
                     32377 => "01011100",
                     32378 => "01010100",
                     32379 => "01001100",
                     32380 => "01011100",
                     32381 => "00011100",
                     32382 => "00011100",
                     32383 => "01011100",
                     32384 => "01011100",
                     32385 => "01011100",
                     32386 => "01011100",
                     32387 => "01011110",
                     32388 => "01010110",
                     32389 => "01001110",
                     32390 => "01011110",
                     32391 => "01010110",
                     32392 => "01001110",
                     32393 => "01011110",
                     32394 => "00011110",
                     32395 => "00011110",
                     32396 => "01011110",
                     32397 => "01011110",
                     32398 => "01011110",
                     32399 => "01011110",
                     32400 => "01100010",
                     32401 => "01011010",
                     32402 => "01010000",
                     32403 => "01100010",
                     32404 => "01011010",
                     32405 => "01010000",
                     32406 => "01100010",
                     32407 => "00100010",
                     32408 => "00100010",
                     32409 => "01100010",
                     32410 => "11100111",
                     32411 => "11100111",
                     32412 => "11100111",
                     32413 => "00101011",
                     32414 => "10000110",
                     32415 => "00010100",
                     32416 => "10000001",
                     32417 => "00010100",
                     32418 => "10000000",
                     32419 => "00010100",
                     32420 => "00010100",
                     32421 => "10000001",
                     32422 => "00010100",
                     32423 => "00010100",
                     32424 => "00010100",
                     32425 => "00010100",
                     32426 => "10000110",
                     32427 => "00010110",
                     32428 => "10000001",
                     32429 => "00010110",
                     32430 => "10000000",
                     32431 => "00010110",
                     32432 => "00010110",
                     32433 => "10000001",
                     32434 => "00010110",
                     32435 => "00010110",
                     32436 => "00010110",
                     32437 => "00010110",
                     32438 => "10000001",
                     32439 => "00101000",
                     32440 => "00100010",
                     32441 => "00011010",
                     32442 => "00101000",
                     32443 => "00100010",
                     32444 => "00011010",
                     32445 => "00101000",
                     32446 => "10000000",
                     32447 => "00101000",
                     32448 => "00101000",
                     32449 => "10000001",
                     32450 => "00101000",
                     32451 => "10000111",
                     32452 => "00101100",
                     32453 => "00101100",
                     32454 => "00101100",
                     32455 => "10000100",
                     32456 => "00110000",
                     32457 => "10000011",
                     32458 => "00000100",
                     32459 => "10000100",
                     32460 => "00001100",
                     32461 => "10000011",
                     32462 => "01100010",
                     32463 => "00010000",
                     32464 => "10000100",
                     32465 => "00010010",
                     32466 => "10000011",
                     32467 => "00011100",
                     32468 => "00100010",
                     32469 => "00011110",
                     32470 => "00100010",
                     32471 => "00100110",
                     32472 => "00011000",
                     32473 => "00011110",
                     32474 => "00000100",
                     32475 => "00011100",
                     32476 => "00000000",
                     32477 => "11100011",
                     32478 => "11100001",
                     32479 => "11100011",
                     32480 => "00011101",
                     32481 => "11011110",
                     32482 => "11100000",
                     32483 => "00100011",
                     32484 => "11101100",
                     32485 => "01110101",
                     32486 => "01110100",
                     32487 => "11110000",
                     32488 => "11110100",
                     32489 => "11110110",
                     32490 => "11101010",
                     32491 => "00110001",
                     32492 => "00101101",
                     32493 => "10000011",
                     32494 => "00010010",
                     32495 => "00010100",
                     32496 => "00000100",
                     32497 => "00011000",
                     32498 => "00011010",
                     32499 => "00011100",
                     32500 => "00010100",
                     32501 => "00100110",
                     32502 => "00100010",
                     32503 => "00011110",
                     32504 => "00011100",
                     32505 => "00011000",
                     32506 => "00011110",
                     32507 => "00100010",
                     32508 => "00001100",
                     32509 => "00010100",
                     32510 => "11111111",
                     32511 => "11111111",
                     32512 => "00000000",
                     32513 => "10001000",
                     32514 => "00000000",
                     32515 => "00101011",
                     32516 => "00000000",
                     32517 => "00000000",
                     32518 => "00000010",
                     32519 => "01110010",
                     32520 => "00000010",
                     32521 => "01001111",
                     32522 => "00000010",
                     32523 => "00101110",
                     32524 => "00000010",
                     32525 => "00001110",
                     32526 => "00000001",
                     32527 => "11110001",
                     32528 => "00000001",
                     32529 => "10111010",
                     32530 => "00000001",
                     32531 => "10100001",
                     32532 => "00000001",
                     32533 => "10001010",
                     32534 => "00000001",
                     32535 => "01110100",
                     32536 => "00000001",
                     32537 => "01011111",
                     32538 => "00000001",
                     32539 => "01001011",
                     32540 => "00000001",
                     32541 => "00111001",
                     32542 => "00000001",
                     32543 => "00100111",
                     32544 => "00000001",
                     32545 => "00010111",
                     32546 => "00000001",
                     32547 => "00000111",
                     32548 => "00000000",
                     32549 => "11111000",
                     32550 => "00000000",
                     32551 => "11101010",
                     32552 => "00000000",
                     32553 => "11011101",
                     32554 => "00000000",
                     32555 => "11010001",
                     32556 => "00000000",
                     32557 => "11000101",
                     32558 => "00000000",
                     32559 => "10111010",
                     32560 => "00000000",
                     32561 => "10101111",
                     32562 => "00000000",
                     32563 => "10100101",
                     32564 => "00000000",
                     32565 => "10011100",
                     32566 => "00000000",
                     32567 => "10010100",
                     32568 => "00000000",
                     32569 => "10001011",
                     32570 => "00000000",
                     32571 => "10000011",
                     32572 => "00000000",
                     32573 => "01111100",
                     32574 => "00000000",
                     32575 => "01101110",
                     32576 => "00000000",
                     32577 => "01110100",
                     32578 => "00000000",
                     32579 => "01101000",
                     32580 => "00000000",
                     32581 => "01001110",
                     32582 => "00000000",
                     32583 => "01011100",
                     32584 => "00000000",
                     32585 => "01011000",
                     32586 => "00000000",
                     32587 => "01010010",
                     32588 => "00000000",
                     32589 => "01001010",
                     32590 => "00000000",
                     32591 => "01000010",
                     32592 => "00000000",
                     32593 => "00111110",
                     32594 => "00000000",
                     32595 => "00110110",
                     32596 => "00000000",
                     32597 => "00110001",
                     32598 => "00000000",
                     32599 => "00100111",
                     32600 => "00000000",
                     32601 => "00100000",
                     32602 => "00000100",
                     32603 => "00011101",
                     32604 => "00000011",
                     32605 => "00010101",
                     32606 => "00000010",
                     32607 => "10111110",
                     32608 => "00000010",
                     32609 => "10011000",
                     32610 => "00000001",
                     32611 => "11010101",
                     32612 => "00000000",
                     32613 => "01100010",
                     32614 => "00000100",
                     32615 => "00001000",
                     32616 => "00010000",
                     32617 => "00100000",
                     32618 => "01000000",
                     32619 => "00011000",
                     32620 => "00110000",
                     32621 => "00001100",
                     32622 => "00000011",
                     32623 => "00000110",
                     32624 => "00001100",
                     32625 => "00011000",
                     32626 => "00110000",
                     32627 => "00010010",
                     32628 => "00100100",
                     32629 => "00001000",
                     32630 => "00000011",
                     32631 => "00000110",
                     32632 => "00001100",
                     32633 => "00011000",
                     32634 => "00110000",
                     32635 => "00010010",
                     32636 => "00100100",
                     32637 => "00001000",
                     32638 => "00100100",
                     32639 => "00000010",
                     32640 => "00000110",
                     32641 => "00000100",
                     32642 => "00001100",
                     32643 => "00010010",
                     32644 => "00011000",
                     32645 => "00001000",
                     32646 => "00011011",
                     32647 => "00000001",
                     32648 => "00000101",
                     32649 => "00000011",
                     32650 => "00001001",
                     32651 => "00001101",
                     32652 => "00010010",
                     32653 => "00000110",
                     32654 => "00010010",
                     32655 => "00000001",
                     32656 => "00000011",
                     32657 => "00000010",
                     32658 => "00000110",
                     32659 => "00001001",
                     32660 => "00001100",
                     32661 => "00000100",
                     32662 => "10011000",
                     32663 => "10011001",
                     32664 => "10011010",
                     32665 => "10011011",
                     32666 => "10010000",
                     32667 => "10010100",
                     32668 => "10010100",
                     32669 => "10010101",
                     32670 => "10010101",
                     32671 => "10010110",
                     32672 => "10010111",
                     32673 => "10011000",
                     32674 => "10010000",
                     32675 => "10010001",
                     32676 => "10010010",
                     32677 => "10010010",
                     32678 => "10010011",
                     32679 => "10010011",
                     32680 => "10010011",
                     32681 => "10010100",
                     32682 => "10010100",
                     32683 => "10010100",
                     32684 => "10010100",
                     32685 => "10010100",
                     32686 => "10010100",
                     32687 => "10010101",
                     32688 => "10010101",
                     32689 => "10010101",
                     32690 => "10010101",
                     32691 => "10010101",
                     32692 => "10010101",
                     32693 => "10010110",
                     32694 => "10010110",
                     32695 => "10010110",
                     32696 => "10010110",
                     32697 => "10010110",
                     32698 => "10010110",
                     32699 => "10010110",
                     32700 => "10010110",
                     32701 => "10010110",
                     32702 => "10010110",
                     32703 => "10010110",
                     32704 => "10010110",
                     32705 => "10010110",
                     32706 => "10010110",
                     32707 => "10010110",
                     32708 => "10010110",
                     32709 => "10010110",
                     32710 => "10010101",
                     32711 => "10010101",
                     32712 => "10010100",
                     32713 => "10010011",
                     32714 => "00010101",
                     32715 => "00010110",
                     32716 => "00010110",
                     32717 => "00010111",
                     32718 => "00010111",
                     32719 => "00011000",
                     32720 => "00011001",
                     32721 => "00011001",
                     32722 => "00011010",
                     32723 => "00011010",
                     32724 => "00011100",
                     32725 => "00011101",
                     32726 => "00011101",
                     32727 => "00011110",
                     32728 => "00011110",
                     32729 => "00011111",
                     32730 => "00011111",
                     32731 => "00011111",
                     32732 => "00011111",
                     32733 => "00011110",
                     32734 => "00011101",
                     32735 => "00011100",
                     32736 => "00011110",
                     32737 => "00011111",
                     32738 => "00011111",
                     32739 => "00011110",
                     32740 => "00011101",
                     32741 => "00011100",
                     32742 => "00011010",
                     32743 => "00011000",
                     32744 => "00010110",
                     32745 => "00010100",
                     32746 => "00010101",
                     32747 => "00010110",
                     32748 => "00010110",
                     32749 => "00010111",
                     32750 => "00010111",
                     32751 => "00011000",
                     32752 => "00011001",
                     32753 => "00011001",
                     32754 => "00011010",
                     32755 => "00011010",
                     32756 => "00011100",
                     32757 => "00011101",
                     32758 => "00011101",
                     32759 => "00011110",
                     32760 => "00011110",
                     32761 => "00011111",
                     32762 => "10000010",
                     32763 => "10000000",
                     32764 => "00000000",
                     32765 => "10000000",
                     32766 => "11110000",
                     32767 => "11111111"
                    );
                                    
                    chr_rom <= (
                     0 => "00000011",
                     1 => "00001111",
                     2 => "00011111",
                     3 => "00011111",
                     4 => "00011100",
                     5 => "00100100",
                     6 => "00100110",
                     7 => "01100110",
                     8 => "00000000",
                     9 => "00000000",
                     10 => "00000000",
                     11 => "00000000",
                     12 => "00011111",
                     13 => "00111111",
                     14 => "00111111",
                     15 => "01111111",
                     16 => "11100000",
                     17 => "11000000",
                     18 => "10000000",
                     19 => "11111100",
                     20 => "10000000",
                     21 => "11000000",
                     22 => "00000000",
                     23 => "00100000",
                     24 => "00000000",
                     25 => "00100000",
                     26 => "01100000",
                     27 => "00000000",
                     28 => "11110000",
                     29 => "11111100",
                     30 => "11111110",
                     31 => "11111110",
                     32 => "01100000",
                     33 => "01110000",
                     34 => "00011000",
                     35 => "00000111",
                     36 => "00001111",
                     37 => "00011111",
                     38 => "00111111",
                     39 => "01111111",
                     40 => "01111111",
                     41 => "01111111",
                     42 => "00011111",
                     43 => "00000111",
                     44 => "00000000",
                     45 => "00011110",
                     46 => "00111111",
                     47 => "01111111",
                     48 => "11111100",
                     49 => "01111100",
                     50 => "00000000",
                     51 => "00000000",
                     52 => "11100000",
                     53 => "11110000",
                     54 => "11111000",
                     55 => "11111000",
                     56 => "11111100",
                     57 => "11111100",
                     58 => "11111000",
                     59 => "11000000",
                     60 => "11000010",
                     61 => "01100111",
                     62 => "00101111",
                     63 => "00110111",
                     64 => "01111111",
                     65 => "01111111",
                     66 => "11111111",
                     67 => "11111111",
                     68 => "00000111",
                     69 => "00000111",
                     70 => "00001111",
                     71 => "00001111",
                     72 => "01111111",
                     73 => "01111110",
                     74 => "11111100",
                     75 => "11110000",
                     76 => "11111000",
                     77 => "11111000",
                     78 => "11110000",
                     79 => "01110000",
                     80 => "11111101",
                     81 => "11111110",
                     82 => "10110100",
                     83 => "11111000",
                     84 => "11111000",
                     85 => "11111001",
                     86 => "11111011",
                     87 => "11111111",
                     88 => "00110111",
                     89 => "00110110",
                     90 => "01011100",
                     91 => "00000000",
                     92 => "00000000",
                     93 => "00000001",
                     94 => "00000011",
                     95 => "00011111",
                     96 => "00011111",
                     97 => "00111111",
                     98 => "11111111",
                     99 => "11111111",
                     100 => "11111100",
                     101 => "01110000",
                     102 => "01110000",
                     103 => "00111000",
                     104 => "00001000",
                     105 => "00100100",
                     106 => "11100011",
                     107 => "11110000",
                     108 => "11111000",
                     109 => "01110000",
                     110 => "01110000",
                     111 => "00111000",
                     112 => "11111111",
                     113 => "11111111",
                     114 => "11111111",
                     115 => "00011111",
                     116 => "00000000",
                     117 => "00000000",
                     118 => "00000000",
                     119 => "00000000",
                     120 => "00011111",
                     121 => "00011111",
                     122 => "00011111",
                     123 => "00011111",
                     124 => "00000000",
                     125 => "00000000",
                     126 => "00000000",
                     127 => "00000000",
                     128 => "00000000",
                     129 => "00000000",
                     130 => "00000001",
                     131 => "00000111",
                     132 => "00001111",
                     133 => "00001111",
                     134 => "00001110",
                     135 => "00010010",
                     136 => "00000000",
                     137 => "00000000",
                     138 => "00000000",
                     139 => "00000000",
                     140 => "00000000",
                     141 => "00000000",
                     142 => "00001111",
                     143 => "00011111",
                     144 => "00000000",
                     145 => "00000000",
                     146 => "11110000",
                     147 => "11100000",
                     148 => "11000000",
                     149 => "11111110",
                     150 => "01000000",
                     151 => "01100000",
                     152 => "00000000",
                     153 => "00000000",
                     154 => "00000000",
                     155 => "00010000",
                     156 => "00110000",
                     157 => "00000000",
                     158 => "11111000",
                     159 => "11111110",
                     160 => "00010011",
                     161 => "00110011",
                     162 => "00110000",
                     163 => "00011000",
                     164 => "00000100",
                     165 => "00001111",
                     166 => "00011111",
                     167 => "00011111",
                     168 => "00011111",
                     169 => "00111111",
                     170 => "00111111",
                     171 => "00011111",
                     172 => "00000111",
                     173 => "00001000",
                     174 => "00010111",
                     175 => "00010111",
                     176 => "00000000",
                     177 => "00010000",
                     178 => "01111110",
                     179 => "00111110",
                     180 => "00000000",
                     181 => "00000000",
                     182 => "11000000",
                     183 => "11100000",
                     184 => "11111111",
                     185 => "11111111",
                     186 => "11111110",
                     187 => "11111110",
                     188 => "11111100",
                     189 => "11100000",
                     190 => "01000000",
                     191 => "10100000",
                     192 => "00111111",
                     193 => "00111111",
                     194 => "00111111",
                     195 => "00011111",
                     196 => "00011111",
                     197 => "00011111",
                     198 => "00011111",
                     199 => "00011111",
                     200 => "00110111",
                     201 => "00100111",
                     202 => "00100011",
                     203 => "00000011",
                     204 => "00000001",
                     205 => "00000000",
                     206 => "00000000",
                     207 => "00000000",
                     208 => "11110000",
                     209 => "11110000",
                     210 => "11110000",
                     211 => "11111000",
                     212 => "11111000",
                     213 => "11111000",
                     214 => "11111000",
                     215 => "11111000",
                     216 => "11001100",
                     217 => "11111111",
                     218 => "11111111",
                     219 => "11111111",
                     220 => "11111111",
                     221 => "01110000",
                     222 => "00000000",
                     223 => "00001000",
                     224 => "11111111",
                     225 => "11111111",
                     226 => "11111111",
                     227 => "11111110",
                     228 => "11110000",
                     229 => "11000000",
                     230 => "10000000",
                     231 => "00000000",
                     232 => "11110000",
                     233 => "11110000",
                     234 => "11110000",
                     235 => "11110000",
                     236 => "11110000",
                     237 => "11000000",
                     238 => "10000000",
                     239 => "00000000",
                     240 => "11111100",
                     241 => "11111100",
                     242 => "11111000",
                     243 => "01111000",
                     244 => "01111000",
                     245 => "01111000",
                     246 => "01111110",
                     247 => "01111110",
                     248 => "00010000",
                     249 => "01100000",
                     250 => "10000000",
                     251 => "00000000",
                     252 => "01111000",
                     253 => "01111000",
                     254 => "01111110",
                     255 => "01111110",
                     256 => "00000000",
                     257 => "00000011",
                     258 => "00001111",
                     259 => "00011111",
                     260 => "00011111",
                     261 => "00011100",
                     262 => "00100100",
                     263 => "00100110",
                     264 => "00000000",
                     265 => "00000000",
                     266 => "00000000",
                     267 => "00000000",
                     268 => "00000000",
                     269 => "00011111",
                     270 => "00111111",
                     271 => "00111111",
                     272 => "00000000",
                     273 => "11100000",
                     274 => "11000000",
                     275 => "10000000",
                     276 => "11111100",
                     277 => "10000000",
                     278 => "11000000",
                     279 => "00000000",
                     280 => "00000000",
                     281 => "00000000",
                     282 => "00100000",
                     283 => "01100000",
                     284 => "00000000",
                     285 => "11110000",
                     286 => "11111100",
                     287 => "11111110",
                     288 => "01100110",
                     289 => "01100000",
                     290 => "00110000",
                     291 => "00011000",
                     292 => "00001111",
                     293 => "00011111",
                     294 => "00111111",
                     295 => "00111111",
                     296 => "01111111",
                     297 => "01111111",
                     298 => "00111111",
                     299 => "00011111",
                     300 => "00000000",
                     301 => "00010110",
                     302 => "00101111",
                     303 => "00101111",
                     304 => "00100000",
                     305 => "11111100",
                     306 => "01111100",
                     307 => "00000000",
                     308 => "00000000",
                     309 => "11100000",
                     310 => "11100000",
                     311 => "11110000",
                     312 => "11111110",
                     313 => "11111100",
                     314 => "11111100",
                     315 => "11111000",
                     316 => "11000000",
                     317 => "01100000",
                     318 => "00100000",
                     319 => "00110000",
                     320 => "00111111",
                     321 => "00111111",
                     322 => "00111111",
                     323 => "00111111",
                     324 => "00111111",
                     325 => "00111111",
                     326 => "00111111",
                     327 => "00011111",
                     328 => "00101111",
                     329 => "00101111",
                     330 => "00101111",
                     331 => "00001111",
                     332 => "00000111",
                     333 => "00000011",
                     334 => "00000000",
                     335 => "00000000",
                     336 => "11110000",
                     337 => "10010000",
                     338 => "00000000",
                     339 => "00001000",
                     340 => "00001100",
                     341 => "00011100",
                     342 => "11111100",
                     343 => "11111000",
                     344 => "00010000",
                     345 => "11110000",
                     346 => "11110000",
                     347 => "11110000",
                     348 => "11110000",
                     349 => "11100000",
                     350 => "11000000",
                     351 => "11100000",
                     352 => "00001111",
                     353 => "00001111",
                     354 => "00000111",
                     355 => "00000111",
                     356 => "00000111",
                     357 => "00001111",
                     358 => "00001111",
                     359 => "00000011",
                     360 => "00000001",
                     361 => "00000011",
                     362 => "00000001",
                     363 => "00000100",
                     364 => "00000111",
                     365 => "00001111",
                     366 => "00001111",
                     367 => "00000011",
                     368 => "11111000",
                     369 => "11110000",
                     370 => "11100000",
                     371 => "11110000",
                     372 => "10110000",
                     373 => "10000000",
                     374 => "11100000",
                     375 => "11100000",
                     376 => "11111000",
                     377 => "11110000",
                     378 => "11100000",
                     379 => "01110000",
                     380 => "10110000",
                     381 => "10000000",
                     382 => "11100000",
                     383 => "11100000",
                     384 => "00000011",
                     385 => "00111111",
                     386 => "01111111",
                     387 => "00011001",
                     388 => "00001001",
                     389 => "00001001",
                     390 => "00101000",
                     391 => "01011100",
                     392 => "00000000",
                     393 => "00110000",
                     394 => "01110000",
                     395 => "01111111",
                     396 => "11111111",
                     397 => "11111111",
                     398 => "11110111",
                     399 => "11110011",
                     400 => "11111000",
                     401 => "11100000",
                     402 => "11100000",
                     403 => "11111100",
                     404 => "00100110",
                     405 => "00110000",
                     406 => "10000000",
                     407 => "00010000",
                     408 => "00000000",
                     409 => "00011000",
                     410 => "00010000",
                     411 => "00000000",
                     412 => "11111000",
                     413 => "11111000",
                     414 => "11111110",
                     415 => "11111111",
                     416 => "00111110",
                     417 => "00011110",
                     418 => "00111111",
                     419 => "00111000",
                     420 => "00110000",
                     421 => "00110000",
                     422 => "00000000",
                     423 => "00111010",
                     424 => "11100111",
                     425 => "00001111",
                     426 => "00001111",
                     427 => "00011111",
                     428 => "00011111",
                     429 => "00011111",
                     430 => "00001111",
                     431 => "00000111",
                     432 => "01111000",
                     433 => "00011110",
                     434 => "10000000",
                     435 => "11111110",
                     436 => "01111110",
                     437 => "01111110",
                     438 => "01111111",
                     439 => "01111111",
                     440 => "11111111",
                     441 => "11111110",
                     442 => "11111100",
                     443 => "11000110",
                     444 => "10001110",
                     445 => "11101110",
                     446 => "11111111",
                     447 => "11111111",
                     448 => "00111100",
                     449 => "00111111",
                     450 => "00011111",
                     451 => "00001111",
                     452 => "00000111",
                     453 => "00111111",
                     454 => "00100001",
                     455 => "00100000",
                     456 => "00000011",
                     457 => "00000000",
                     458 => "00000000",
                     459 => "00001110",
                     460 => "00000111",
                     461 => "00111111",
                     462 => "00111111",
                     463 => "00111111",
                     464 => "11111111",
                     465 => "11111111",
                     466 => "11111111",
                     467 => "11111110",
                     468 => "11111110",
                     469 => "11111110",
                     470 => "11111100",
                     471 => "01110000",
                     472 => "11111111",
                     473 => "01111111",
                     474 => "00111111",
                     475 => "00001110",
                     476 => "11000000",
                     477 => "11000000",
                     478 => "11100000",
                     479 => "11100000",
                     480 => "00001111",
                     481 => "10011111",
                     482 => "11001111",
                     483 => "11111111",
                     484 => "01111111",
                     485 => "00111111",
                     486 => "00011110",
                     487 => "00001110",
                     488 => "00000000",
                     489 => "10000000",
                     490 => "11001000",
                     491 => "11111110",
                     492 => "01111111",
                     493 => "00111111",
                     494 => "00011110",
                     495 => "00001110",
                     496 => "00100000",
                     497 => "11000000",
                     498 => "10000000",
                     499 => "10000000",
                     500 => "00000000",
                     501 => "00000000",
                     502 => "00000000",
                     503 => "00000000",
                     504 => "11100000",
                     505 => "00000000",
                     506 => "00000000",
                     507 => "00000000",
                     508 => "00000000",
                     509 => "00000000",
                     510 => "00000000",
                     511 => "00000000",
                     512 => "00000000",
                     513 => "00000000",
                     514 => "00000011",
                     515 => "00001111",
                     516 => "00011111",
                     517 => "00011111",
                     518 => "00011100",
                     519 => "00100100",
                     520 => "00000000",
                     521 => "00000000",
                     522 => "00000000",
                     523 => "00000000",
                     524 => "00000000",
                     525 => "00000000",
                     526 => "00011111",
                     527 => "00111111",
                     528 => "00000000",
                     529 => "00000100",
                     530 => "11100110",
                     531 => "11100000",
                     532 => "11111111",
                     533 => "11111111",
                     534 => "10001111",
                     535 => "10000011",
                     536 => "00001110",
                     537 => "00011111",
                     538 => "00011111",
                     539 => "00011111",
                     540 => "00011111",
                     541 => "00000011",
                     542 => "11111111",
                     543 => "11111111",
                     544 => "00100110",
                     545 => "00100110",
                     546 => "01100000",
                     547 => "01111000",
                     548 => "00011000",
                     549 => "00001111",
                     550 => "01111111",
                     551 => "11111111",
                     552 => "00111111",
                     553 => "00111111",
                     554 => "01111111",
                     555 => "01111111",
                     556 => "00011111",
                     557 => "00000000",
                     558 => "01111110",
                     559 => "11111111",
                     560 => "00000001",
                     561 => "00100001",
                     562 => "11111110",
                     563 => "01111010",
                     564 => "00000110",
                     565 => "11111110",
                     566 => "11111100",
                     567 => "11111100",
                     568 => "11111111",
                     569 => "11111111",
                     570 => "11111110",
                     571 => "11111110",
                     572 => "11111110",
                     573 => "11011110",
                     574 => "01011100",
                     575 => "01101100",
                     576 => "11111111",
                     577 => "11001111",
                     578 => "10000111",
                     579 => "00000111",
                     580 => "00000111",
                     581 => "00001111",
                     582 => "00011111",
                     583 => "00011111",
                     584 => "11111111",
                     585 => "11111111",
                     586 => "11111110",
                     587 => "11111100",
                     588 => "11111000",
                     589 => "10110000",
                     590 => "01100000",
                     591 => "00000000",
                     592 => "11111000",
                     593 => "11111000",
                     594 => "11110000",
                     595 => "10111000",
                     596 => "11111000",
                     597 => "11111001",
                     598 => "11111011",
                     599 => "11111111",
                     600 => "00101000",
                     601 => "00110000",
                     602 => "00011000",
                     603 => "01000000",
                     604 => "00000000",
                     605 => "00000001",
                     606 => "00000011",
                     607 => "00001111",
                     608 => "00011111",
                     609 => "11111111",
                     610 => "11111111",
                     611 => "11111111",
                     612 => "11111111",
                     613 => "11111110",
                     614 => "11000000",
                     615 => "10000000",
                     616 => "00010000",
                     617 => "11101100",
                     618 => "11100011",
                     619 => "11100000",
                     620 => "11100000",
                     621 => "11100000",
                     622 => "11000000",
                     623 => "10000000",
                     624 => "11111111",
                     625 => "11111111",
                     626 => "11111111",
                     627 => "00111111",
                     628 => "00000000",
                     629 => "00000000",
                     630 => "00000000",
                     631 => "00000000",
                     632 => "00001111",
                     633 => "00001111",
                     634 => "00001111",
                     635 => "00001111",
                     636 => "00000000",
                     637 => "00000000",
                     638 => "00000000",
                     639 => "00000000",
                     640 => "00010011",
                     641 => "00110011",
                     642 => "00110000",
                     643 => "00011000",
                     644 => "00000100",
                     645 => "00001111",
                     646 => "00011111",
                     647 => "00011111",
                     648 => "00011111",
                     649 => "00111111",
                     650 => "00111111",
                     651 => "00011111",
                     652 => "00000111",
                     653 => "00001001",
                     654 => "00010011",
                     655 => "00010111",
                     656 => "00000000",
                     657 => "00010000",
                     658 => "01111110",
                     659 => "00110000",
                     660 => "11100000",
                     661 => "11110000",
                     662 => "11110000",
                     663 => "11100000",
                     664 => "11111111",
                     665 => "11111111",
                     666 => "11111110",
                     667 => "11111111",
                     668 => "11111110",
                     669 => "11111100",
                     670 => "11111000",
                     671 => "11100000",
                     672 => "00011111",
                     673 => "00011111",
                     674 => "00001111",
                     675 => "00001111",
                     676 => "00001111",
                     677 => "00011111",
                     678 => "00011111",
                     679 => "00011111",
                     680 => "00010111",
                     681 => "00010111",
                     682 => "00000011",
                     683 => "00000000",
                     684 => "00000000",
                     685 => "00000000",
                     686 => "00000000",
                     687 => "00000000",
                     688 => "11110000",
                     689 => "11110000",
                     690 => "11111000",
                     691 => "11111000",
                     692 => "10111000",
                     693 => "11111000",
                     694 => "11111000",
                     695 => "11111000",
                     696 => "11010000",
                     697 => "10010000",
                     698 => "00011000",
                     699 => "00001000",
                     700 => "01000000",
                     701 => "00000000",
                     702 => "00000000",
                     703 => "00000000",
                     704 => "00111111",
                     705 => "11111111",
                     706 => "11111111",
                     707 => "11111111",
                     708 => "11110110",
                     709 => "11000110",
                     710 => "10000100",
                     711 => "00000000",
                     712 => "00110000",
                     713 => "11110000",
                     714 => "11110000",
                     715 => "11110001",
                     716 => "11110110",
                     717 => "11000110",
                     718 => "10000100",
                     719 => "00000000",
                     720 => "11110000",
                     721 => "11100000",
                     722 => "10000000",
                     723 => "00000000",
                     724 => "00000000",
                     725 => "00000000",
                     726 => "00000000",
                     727 => "00000000",
                     728 => "00000000",
                     729 => "00000000",
                     730 => "00000000",
                     731 => "00000000",
                     732 => "00000000",
                     733 => "00000000",
                     734 => "00000000",
                     735 => "00000000",
                     736 => "00011111",
                     737 => "00011111",
                     738 => "00111111",
                     739 => "00111111",
                     740 => "00011111",
                     741 => "00001111",
                     742 => "00001111",
                     743 => "00011111",
                     744 => "00011111",
                     745 => "00011111",
                     746 => "00111111",
                     747 => "00111110",
                     748 => "01111100",
                     749 => "01111000",
                     750 => "11110000",
                     751 => "11100000",
                     752 => "11110000",
                     753 => "11110000",
                     754 => "11111000",
                     755 => "11111000",
                     756 => "10111000",
                     757 => "11111000",
                     758 => "11111000",
                     759 => "11110000",
                     760 => "10110000",
                     761 => "10010000",
                     762 => "00011000",
                     763 => "00001000",
                     764 => "01000000",
                     765 => "00000000",
                     766 => "00000000",
                     767 => "00000000",
                     768 => "11100000",
                     769 => "11110000",
                     770 => "11110000",
                     771 => "11110000",
                     772 => "11110000",
                     773 => "11110000",
                     774 => "11111000",
                     775 => "11110000",
                     776 => "11000000",
                     777 => "11100000",
                     778 => "11111100",
                     779 => "11111110",
                     780 => "11111111",
                     781 => "01111111",
                     782 => "00000011",
                     783 => "00000000",
                     784 => "00011111",
                     785 => "00011111",
                     786 => "00011111",
                     787 => "00111111",
                     788 => "00111110",
                     789 => "00111100",
                     790 => "00111000",
                     791 => "00011000",
                     792 => "00000000",
                     793 => "00000000",
                     794 => "00010000",
                     795 => "00111000",
                     796 => "00111110",
                     797 => "00111100",
                     798 => "00111000",
                     799 => "00011000",
                     800 => "00000000",
                     801 => "00000011",
                     802 => "00000111",
                     803 => "00000111",
                     804 => "00001010",
                     805 => "00001011",
                     806 => "00001100",
                     807 => "00000000",
                     808 => "00000000",
                     809 => "00000000",
                     810 => "00000000",
                     811 => "00000111",
                     812 => "00001111",
                     813 => "00001111",
                     814 => "00001111",
                     815 => "00000011",
                     816 => "00000000",
                     817 => "11100000",
                     818 => "11111100",
                     819 => "00100000",
                     820 => "00100000",
                     821 => "00010000",
                     822 => "00111100",
                     823 => "00000000",
                     824 => "00000000",
                     825 => "00000000",
                     826 => "00000000",
                     827 => "11110000",
                     828 => "11111100",
                     829 => "11111110",
                     830 => "11111100",
                     831 => "11111000",
                     832 => "00000111",
                     833 => "00000111",
                     834 => "00000111",
                     835 => "00011111",
                     836 => "00011111",
                     837 => "00111110",
                     838 => "00100001",
                     839 => "00000001",
                     840 => "00000111",
                     841 => "00001111",
                     842 => "00011011",
                     843 => "00011000",
                     844 => "00010000",
                     845 => "00110000",
                     846 => "00100001",
                     847 => "00000001",
                     848 => "11100000",
                     849 => "11100000",
                     850 => "11100000",
                     851 => "11110000",
                     852 => "11110000",
                     853 => "11100000",
                     854 => "11000000",
                     855 => "11100000",
                     856 => "10101000",
                     857 => "11111100",
                     858 => "11111000",
                     859 => "00000000",
                     860 => "00000000",
                     861 => "00000000",
                     862 => "11000000",
                     863 => "11100000",
                     864 => "00000111",
                     865 => "00001111",
                     866 => "00001110",
                     867 => "00010100",
                     868 => "00010110",
                     869 => "00011000",
                     870 => "00000000",
                     871 => "00111111",
                     872 => "00000000",
                     873 => "00000000",
                     874 => "00001111",
                     875 => "00011111",
                     876 => "00011111",
                     877 => "00011111",
                     878 => "00000111",
                     879 => "00111100",
                     880 => "11000000",
                     881 => "11111000",
                     882 => "01000000",
                     883 => "01000000",
                     884 => "00100000",
                     885 => "01111000",
                     886 => "00000000",
                     887 => "11000000",
                     888 => "00000000",
                     889 => "00000000",
                     890 => "11100000",
                     891 => "11111000",
                     892 => "11111100",
                     893 => "11111000",
                     894 => "11110000",
                     895 => "11000000",
                     896 => "00111111",
                     897 => "00001110",
                     898 => "00001111",
                     899 => "00011111",
                     900 => "00111111",
                     901 => "01111100",
                     902 => "01110000",
                     903 => "00111000",
                     904 => "11111100",
                     905 => "11101101",
                     906 => "11000000",
                     907 => "00000000",
                     908 => "00000000",
                     909 => "01100000",
                     910 => "01110000",
                     911 => "00111000",
                     912 => "11110000",
                     913 => "11111000",
                     914 => "11100100",
                     915 => "11111100",
                     916 => "11111100",
                     917 => "01111100",
                     918 => "00000000",
                     919 => "00000000",
                     920 => "01111110",
                     921 => "00011110",
                     922 => "00000100",
                     923 => "00001100",
                     924 => "00001100",
                     925 => "00001100",
                     926 => "00000000",
                     927 => "00000000",
                     928 => "00000111",
                     929 => "00001111",
                     930 => "00001110",
                     931 => "00010100",
                     932 => "00010110",
                     933 => "00011000",
                     934 => "00000000",
                     935 => "00001111",
                     936 => "00000000",
                     937 => "00000000",
                     938 => "00001111",
                     939 => "00011111",
                     940 => "00011111",
                     941 => "00011111",
                     942 => "00000111",
                     943 => "00001101",
                     944 => "00011111",
                     945 => "00011111",
                     946 => "00011111",
                     947 => "00011100",
                     948 => "00001100",
                     949 => "00000111",
                     950 => "00000111",
                     951 => "00000111",
                     952 => "00011110",
                     953 => "00011100",
                     954 => "00011110",
                     955 => "00001111",
                     956 => "00000111",
                     957 => "00000000",
                     958 => "00000111",
                     959 => "00000111",
                     960 => "11100000",
                     961 => "01100000",
                     962 => "11110000",
                     963 => "01110000",
                     964 => "11100000",
                     965 => "11100000",
                     966 => "11110000",
                     967 => "10000000",
                     968 => "01100000",
                     969 => "10010000",
                     970 => "00000000",
                     971 => "10000000",
                     972 => "00000000",
                     973 => "11100000",
                     974 => "11110000",
                     975 => "10000000",
                     976 => "00000111",
                     977 => "00011111",
                     978 => "00111111",
                     979 => "00010010",
                     980 => "00010011",
                     981 => "00001000",
                     982 => "00011111",
                     983 => "00110001",
                     984 => "00000000",
                     985 => "00010000",
                     986 => "00111111",
                     987 => "01111111",
                     988 => "01111111",
                     989 => "00111111",
                     990 => "00000011",
                     991 => "00001111",
                     992 => "11000000",
                     993 => "11110000",
                     994 => "01000000",
                     995 => "00000000",
                     996 => "00110000",
                     997 => "00011000",
                     998 => "11000000",
                     999 => "11111000",
                     1000 => "00000000",
                     1001 => "00000000",
                     1002 => "11100000",
                     1003 => "11111000",
                     1004 => "11111100",
                     1005 => "11111000",
                     1006 => "10110000",
                     1007 => "00111000",
                     1008 => "00110001",
                     1009 => "00111001",
                     1010 => "00011111",
                     1011 => "00011111",
                     1012 => "00001111",
                     1013 => "01011111",
                     1014 => "01111110",
                     1015 => "00111100",
                     1016 => "00011111",
                     1017 => "00000111",
                     1018 => "00000000",
                     1019 => "00001110",
                     1020 => "00001111",
                     1021 => "01010011",
                     1022 => "01111100",
                     1023 => "00111100",
                     1024 => "11111000",
                     1025 => "11111000",
                     1026 => "11110000",
                     1027 => "11100000",
                     1028 => "11100000",
                     1029 => "11000000",
                     1030 => "00000000",
                     1031 => "00000000",
                     1032 => "11111000",
                     1033 => "11111000",
                     1034 => "11110000",
                     1035 => "00000000",
                     1036 => "00000000",
                     1037 => "10000000",
                     1038 => "00000000",
                     1039 => "00000000",
                     1040 => "00000000",
                     1041 => "11100000",
                     1042 => "11111100",
                     1043 => "00100111",
                     1044 => "00100111",
                     1045 => "00010001",
                     1046 => "00111110",
                     1047 => "00000100",
                     1048 => "00000111",
                     1049 => "00000111",
                     1050 => "00000011",
                     1051 => "11110111",
                     1052 => "11111111",
                     1053 => "11111111",
                     1054 => "11111110",
                     1055 => "11111100",
                     1056 => "00111111",
                     1057 => "01111111",
                     1058 => "00111111",
                     1059 => "00001111",
                     1060 => "00011111",
                     1061 => "00111111",
                     1062 => "01111111",
                     1063 => "01001111",
                     1064 => "00111110",
                     1065 => "01111111",
                     1066 => "11111111",
                     1067 => "11100010",
                     1068 => "01010000",
                     1069 => "00111000",
                     1070 => "01110000",
                     1071 => "01000000",
                     1072 => "11111000",
                     1073 => "11111001",
                     1074 => "11111001",
                     1075 => "10110111",
                     1076 => "11111111",
                     1077 => "11111111",
                     1078 => "11100000",
                     1079 => "00000000",
                     1080 => "11101000",
                     1081 => "01110001",
                     1082 => "00000001",
                     1083 => "01001011",
                     1084 => "00000011",
                     1085 => "00000011",
                     1086 => "00000000",
                     1087 => "00000000",
                     1088 => "00000111",
                     1089 => "00000111",
                     1090 => "00001111",
                     1091 => "00111111",
                     1092 => "00111111",
                     1093 => "00111111",
                     1094 => "00100110",
                     1095 => "00000100",
                     1096 => "00000101",
                     1097 => "00000011",
                     1098 => "00000001",
                     1099 => "00110000",
                     1100 => "00110000",
                     1101 => "00110000",
                     1102 => "00100110",
                     1103 => "00000100",
                     1104 => "11110000",
                     1105 => "11110000",
                     1106 => "11110000",
                     1107 => "11100000",
                     1108 => "11000000",
                     1109 => "00000000",
                     1110 => "00000000",
                     1111 => "00000000",
                     1112 => "11111110",
                     1113 => "11111100",
                     1114 => "11100000",
                     1115 => "00000000",
                     1116 => "00000000",
                     1117 => "00000000",
                     1118 => "00000000",
                     1119 => "00000000",
                     1120 => "00000111",
                     1121 => "00000111",
                     1122 => "00001111",
                     1123 => "00011111",
                     1124 => "00111111",
                     1125 => "00001111",
                     1126 => "00011100",
                     1127 => "00011000",
                     1128 => "00000101",
                     1129 => "00000011",
                     1130 => "00000001",
                     1131 => "00010000",
                     1132 => "00110000",
                     1133 => "00001100",
                     1134 => "00011100",
                     1135 => "00011000",
                     1136 => "11100000",
                     1137 => "11100000",
                     1138 => "11100000",
                     1139 => "11100000",
                     1140 => "11000000",
                     1141 => "10000000",
                     1142 => "00000000",
                     1143 => "00000000",
                     1144 => "11000000",
                     1145 => "11100000",
                     1146 => "11110000",
                     1147 => "01111000",
                     1148 => "00011000",
                     1149 => "00001000",
                     1150 => "00000000",
                     1151 => "00000000",
                     1152 => "00000111",
                     1153 => "00001111",
                     1154 => "00011111",
                     1155 => "00001111",
                     1156 => "00111111",
                     1157 => "00001111",
                     1158 => "00011100",
                     1159 => "00011000",
                     1160 => "00000111",
                     1161 => "00001111",
                     1162 => "00111110",
                     1163 => "01111100",
                     1164 => "00110000",
                     1165 => "00001100",
                     1166 => "00011100",
                     1167 => "00011000",
                     1168 => "11100000",
                     1169 => "11100000",
                     1170 => "11100000",
                     1171 => "01000000",
                     1172 => "11000000",
                     1173 => "10000000",
                     1174 => "00000000",
                     1175 => "00000000",
                     1176 => "01100000",
                     1177 => "01100000",
                     1178 => "01100000",
                     1179 => "10000000",
                     1180 => "00000000",
                     1181 => "00000000",
                     1182 => "00000000",
                     1183 => "00000000",
                     1184 => "01111111",
                     1185 => "11111111",
                     1186 => "11111111",
                     1187 => "11111011",
                     1188 => "00001111",
                     1189 => "00001111",
                     1190 => "00001111",
                     1191 => "00011111",
                     1192 => "01110011",
                     1193 => "11110011",
                     1194 => "11110000",
                     1195 => "11110100",
                     1196 => "11110000",
                     1197 => "11110000",
                     1198 => "01110000",
                     1199 => "01100000",
                     1200 => "00111111",
                     1201 => "01111110",
                     1202 => "01111100",
                     1203 => "01111100",
                     1204 => "00111100",
                     1205 => "00111100",
                     1206 => "11111100",
                     1207 => "11111100",
                     1208 => "00000000",
                     1209 => "00000000",
                     1210 => "00000000",
                     1211 => "00000000",
                     1212 => "00111100",
                     1213 => "00111100",
                     1214 => "11111100",
                     1215 => "11111100",
                     1216 => "01100000",
                     1217 => "01110000",
                     1218 => "00011000",
                     1219 => "00001000",
                     1220 => "00001111",
                     1221 => "00011111",
                     1222 => "00111111",
                     1223 => "01111111",
                     1224 => "01111111",
                     1225 => "01111111",
                     1226 => "00011111",
                     1227 => "00000111",
                     1228 => "00001011",
                     1229 => "00011011",
                     1230 => "00111011",
                     1231 => "01111011",
                     1232 => "11111100",
                     1233 => "01111100",
                     1234 => "00000000",
                     1235 => "00100000",
                     1236 => "11110000",
                     1237 => "11111000",
                     1238 => "11111100",
                     1239 => "11111110",
                     1240 => "11111100",
                     1241 => "11111100",
                     1242 => "11111000",
                     1243 => "11100000",
                     1244 => "11010000",
                     1245 => "11011000",
                     1246 => "11011100",
                     1247 => "11011110",
                     1248 => "00001011",
                     1249 => "00001111",
                     1250 => "00011111",
                     1251 => "00011110",
                     1252 => "00111100",
                     1253 => "00111100",
                     1254 => "00111100",
                     1255 => "01111100",
                     1256 => "11000100",
                     1257 => "11100000",
                     1258 => "11100000",
                     1259 => "01000000",
                     1260 => "00000000",
                     1261 => "00111100",
                     1262 => "00111100",
                     1263 => "01111100",
                     1264 => "00011111",
                     1265 => "00111111",
                     1266 => "00001101",
                     1267 => "00000111",
                     1268 => "00001111",
                     1269 => "00001110",
                     1270 => "00011100",
                     1271 => "00111100",
                     1272 => "00011101",
                     1273 => "00111100",
                     1274 => "00111010",
                     1275 => "00111000",
                     1276 => "00110000",
                     1277 => "00000000",
                     1278 => "00011100",
                     1279 => "00111100",
                     1280 => "00000000",
                     1281 => "00000000",
                     1282 => "00000000",
                     1283 => "00000000",
                     1284 => "00000000",
                     1285 => "00000000",
                     1286 => "00000000",
                     1287 => "00000000",
                     1288 => "00100010",
                     1289 => "01010101",
                     1290 => "01010101",
                     1291 => "01010101",
                     1292 => "01010101",
                     1293 => "01010101",
                     1294 => "01110111",
                     1295 => "00100010",
                     1296 => "00000000",
                     1297 => "00000111",
                     1298 => "00011111",
                     1299 => "11111111",
                     1300 => "00000111",
                     1301 => "00011111",
                     1302 => "00001111",
                     1303 => "00000110",
                     1304 => "00000000",
                     1305 => "00000000",
                     1306 => "00000000",
                     1307 => "00000000",
                     1308 => "00000000",
                     1309 => "00000000",
                     1310 => "00000000",
                     1311 => "00000000",
                     1312 => "00111111",
                     1313 => "11111111",
                     1314 => "11111111",
                     1315 => "11111111",
                     1316 => "11111111",
                     1317 => "11111111",
                     1318 => "11111011",
                     1319 => "01110110",
                     1320 => "00000000",
                     1321 => "00000000",
                     1322 => "11001111",
                     1323 => "00000111",
                     1324 => "01111111",
                     1325 => "00000000",
                     1326 => "00000000",
                     1327 => "00000000",
                     1328 => "00100000",
                     1329 => "11111000",
                     1330 => "11111111",
                     1331 => "11000011",
                     1332 => "11111101",
                     1333 => "11111110",
                     1334 => "11110000",
                     1335 => "01000000",
                     1336 => "00000000",
                     1337 => "00000000",
                     1338 => "00111100",
                     1339 => "11111100",
                     1340 => "11111110",
                     1341 => "11100000",
                     1342 => "00000000",
                     1343 => "00000000",
                     1344 => "01000000",
                     1345 => "11100000",
                     1346 => "01000000",
                     1347 => "01000000",
                     1348 => "01000001",
                     1349 => "01000001",
                     1350 => "01001111",
                     1351 => "01000111",
                     1352 => "01000000",
                     1353 => "11100000",
                     1354 => "01000000",
                     1355 => "00111111",
                     1356 => "00111110",
                     1357 => "00111110",
                     1358 => "00110000",
                     1359 => "00111000",
                     1360 => "00000000",
                     1361 => "00000000",
                     1362 => "00000000",
                     1363 => "00000000",
                     1364 => "00000000",
                     1365 => "00000000",
                     1366 => "11100000",
                     1367 => "11000000",
                     1368 => "00000000",
                     1369 => "00000000",
                     1370 => "00000000",
                     1371 => "11111000",
                     1372 => "11111000",
                     1373 => "11111000",
                     1374 => "00011000",
                     1375 => "00111000",
                     1376 => "01000011",
                     1377 => "01000110",
                     1378 => "01000100",
                     1379 => "01000000",
                     1380 => "01000000",
                     1381 => "01000000",
                     1382 => "01000000",
                     1383 => "01000000",
                     1384 => "00111100",
                     1385 => "00111001",
                     1386 => "00111011",
                     1387 => "00111111",
                     1388 => "00000000",
                     1389 => "00000000",
                     1390 => "00000000",
                     1391 => "00000000",
                     1392 => "10000000",
                     1393 => "11000000",
                     1394 => "01000000",
                     1395 => "00000000",
                     1396 => "00000000",
                     1397 => "00000000",
                     1398 => "00000000",
                     1399 => "00000000",
                     1400 => "01111000",
                     1401 => "00111000",
                     1402 => "10111000",
                     1403 => "11111000",
                     1404 => "00000000",
                     1405 => "00000000",
                     1406 => "00000000",
                     1407 => "00000000",
                     1408 => "00110001",
                     1409 => "00110000",
                     1410 => "00111000",
                     1411 => "01111100",
                     1412 => "01111111",
                     1413 => "11111111",
                     1414 => "11111111",
                     1415 => "11111011",
                     1416 => "00111111",
                     1417 => "00111111",
                     1418 => "00001111",
                     1419 => "01110111",
                     1420 => "01110111",
                     1421 => "11110111",
                     1422 => "11110111",
                     1423 => "11110111",
                     1424 => "00010000",
                     1425 => "01111110",
                     1426 => "00111110",
                     1427 => "00000000",
                     1428 => "00011110",
                     1429 => "11111110",
                     1430 => "11111111",
                     1431 => "11111111",
                     1432 => "11111111",
                     1433 => "11111110",
                     1434 => "11111110",
                     1435 => "11111110",
                     1436 => "11111010",
                     1437 => "11111010",
                     1438 => "11110011",
                     1439 => "11100111",
                     1440 => "11111111",
                     1441 => "11111111",
                     1442 => "11100011",
                     1443 => "11000011",
                     1444 => "10000111",
                     1445 => "01001000",
                     1446 => "00111100",
                     1447 => "11111100",
                     1448 => "11110000",
                     1449 => "11111000",
                     1450 => "11111100",
                     1451 => "01111100",
                     1452 => "01111000",
                     1453 => "00111000",
                     1454 => "00111100",
                     1455 => "11111100",
                     1456 => "00000000",
                     1457 => "11111111",
                     1458 => "11000011",
                     1459 => "10000011",
                     1460 => "10000011",
                     1461 => "11111111",
                     1462 => "11111111",
                     1463 => "11111111",
                     1464 => "11111111",
                     1465 => "00000000",
                     1466 => "11000011",
                     1467 => "10000001",
                     1468 => "10000001",
                     1469 => "11000011",
                     1470 => "11111111",
                     1471 => "00000000",
                     1472 => "00011111",
                     1473 => "00011111",
                     1474 => "00001111",
                     1475 => "00000111",
                     1476 => "00000001",
                     1477 => "00000000",
                     1478 => "00000000",
                     1479 => "00000000",
                     1480 => "00000000",
                     1481 => "00000000",
                     1482 => "00000000",
                     1483 => "00000000",
                     1484 => "00000000",
                     1485 => "00000000",
                     1486 => "00000000",
                     1487 => "00000000",
                     1488 => "11110000",
                     1489 => "11111011",
                     1490 => "11111111",
                     1491 => "11111111",
                     1492 => "11111110",
                     1493 => "00111110",
                     1494 => "00001100",
                     1495 => "00000100",
                     1496 => "00000000",
                     1497 => "00001011",
                     1498 => "00011111",
                     1499 => "00011111",
                     1500 => "00011110",
                     1501 => "00111110",
                     1502 => "00001100",
                     1503 => "00000100",
                     1504 => "00011111",
                     1505 => "00011111",
                     1506 => "00001111",
                     1507 => "00001111",
                     1508 => "00000111",
                     1509 => "00000000",
                     1510 => "00000000",
                     1511 => "00000000",
                     1512 => "00000000",
                     1513 => "00000000",
                     1514 => "00000000",
                     1515 => "00000000",
                     1516 => "00000000",
                     1517 => "00000000",
                     1518 => "00000000",
                     1519 => "00000000",
                     1520 => "11111011",
                     1521 => "11111111",
                     1522 => "11111111",
                     1523 => "11111111",
                     1524 => "11111111",
                     1525 => "00000000",
                     1526 => "00000000",
                     1527 => "00000000",
                     1528 => "00000011",
                     1529 => "00001111",
                     1530 => "00001111",
                     1531 => "00001111",
                     1532 => "00001111",
                     1533 => "00000000",
                     1534 => "00000000",
                     1535 => "00000000",
                     1536 => "00000000",
                     1537 => "00011000",
                     1538 => "00111100",
                     1539 => "01111110",
                     1540 => "01101110",
                     1541 => "11011111",
                     1542 => "11011111",
                     1543 => "11011111",
                     1544 => "00000000",
                     1545 => "00011000",
                     1546 => "00111100",
                     1547 => "01111110",
                     1548 => "01110110",
                     1549 => "11111011",
                     1550 => "11111011",
                     1551 => "11111011",
                     1552 => "00000000",
                     1553 => "00011000",
                     1554 => "00011000",
                     1555 => "00111100",
                     1556 => "00111100",
                     1557 => "00111100",
                     1558 => "00111100",
                     1559 => "00011100",
                     1560 => "00000000",
                     1561 => "00010000",
                     1562 => "00010000",
                     1563 => "00100000",
                     1564 => "00100000",
                     1565 => "00100000",
                     1566 => "00100000",
                     1567 => "00100000",
                     1568 => "00000000",
                     1569 => "00001000",
                     1570 => "00001000",
                     1571 => "00001000",
                     1572 => "00001000",
                     1573 => "00001000",
                     1574 => "00001000",
                     1575 => "00000000",
                     1576 => "00000000",
                     1577 => "00001000",
                     1578 => "00001000",
                     1579 => "00001000",
                     1580 => "00001000",
                     1581 => "00001000",
                     1582 => "00001000",
                     1583 => "00001000",
                     1584 => "00000000",
                     1585 => "00001000",
                     1586 => "00001000",
                     1587 => "00000100",
                     1588 => "00000100",
                     1589 => "00000100",
                     1590 => "00000100",
                     1591 => "00000100",
                     1592 => "00000000",
                     1593 => "00010000",
                     1594 => "00010000",
                     1595 => "00111000",
                     1596 => "00111000",
                     1597 => "00111000",
                     1598 => "00111000",
                     1599 => "00111000",
                     1600 => "00111100",
                     1601 => "01111110",
                     1602 => "01110111",
                     1603 => "11111011",
                     1604 => "10011111",
                     1605 => "01011111",
                     1606 => "10001110",
                     1607 => "00100000",
                     1608 => "00000000",
                     1609 => "00011000",
                     1610 => "00111100",
                     1611 => "00001110",
                     1612 => "00001110",
                     1613 => "00000100",
                     1614 => "00000000",
                     1615 => "00000000",
                     1616 => "01011100",
                     1617 => "00101110",
                     1618 => "10001111",
                     1619 => "00111111",
                     1620 => "01111011",
                     1621 => "01110111",
                     1622 => "01111110",
                     1623 => "00111100",
                     1624 => "00000000",
                     1625 => "00000000",
                     1626 => "00000100",
                     1627 => "00000110",
                     1628 => "00011110",
                     1629 => "00111100",
                     1630 => "00011000",
                     1631 => "00000000",
                     1632 => "00010011",
                     1633 => "01001111",
                     1634 => "00111111",
                     1635 => "10111111",
                     1636 => "00111111",
                     1637 => "01111010",
                     1638 => "11111000",
                     1639 => "11111000",
                     1640 => "00000000",
                     1641 => "00000000",
                     1642 => "00000001",
                     1643 => "00001010",
                     1644 => "00010111",
                     1645 => "00001111",
                     1646 => "00101111",
                     1647 => "00011111",
                     1648 => "00000000",
                     1649 => "00001000",
                     1650 => "00000101",
                     1651 => "00001111",
                     1652 => "00101111",
                     1653 => "00011101",
                     1654 => "00011100",
                     1655 => "00111100",
                     1656 => "00000000",
                     1657 => "00000000",
                     1658 => "00000000",
                     1659 => "00000000",
                     1660 => "00000101",
                     1661 => "00000111",
                     1662 => "00001111",
                     1663 => "00000111",
                     1664 => "00000000",
                     1665 => "00000000",
                     1666 => "00000000",
                     1667 => "00000000",
                     1668 => "00000010",
                     1669 => "00001011",
                     1670 => "00000111",
                     1671 => "00001111",
                     1672 => "00000000",
                     1673 => "00000000",
                     1674 => "00000000",
                     1675 => "00000000",
                     1676 => "00000000",
                     1677 => "00000000",
                     1678 => "00000001",
                     1679 => "00000011",
                     1680 => "00000000",
                     1681 => "00000000",
                     1682 => "00000000",
                     1683 => "00000000",
                     1684 => "00000000",
                     1685 => "00001000",
                     1686 => "00000100",
                     1687 => "00000100",
                     1688 => "00000000",
                     1689 => "01100000",
                     1690 => "11110000",
                     1691 => "11111000",
                     1692 => "01111100",
                     1693 => "00111110",
                     1694 => "01111110",
                     1695 => "01111111",
                     1696 => "00000010",
                     1697 => "00000010",
                     1698 => "00000010",
                     1699 => "00000101",
                     1700 => "01110001",
                     1701 => "01111111",
                     1702 => "01111111",
                     1703 => "01111111",
                     1704 => "00111111",
                     1705 => "01011111",
                     1706 => "01111111",
                     1707 => "00111110",
                     1708 => "00001110",
                     1709 => "00001010",
                     1710 => "01010001",
                     1711 => "00100000",
                     1712 => "00000000",
                     1713 => "00000000",
                     1714 => "00000000",
                     1715 => "00000000",
                     1716 => "00000000",
                     1717 => "00000000",
                     1718 => "00000000",
                     1719 => "00000100",
                     1720 => "00000000",
                     1721 => "00000000",
                     1722 => "00000000",
                     1723 => "00000000",
                     1724 => "00000000",
                     1725 => "00000000",
                     1726 => "00001110",
                     1727 => "00011111",
                     1728 => "00000010",
                     1729 => "00000010",
                     1730 => "00000000",
                     1731 => "00000001",
                     1732 => "00010011",
                     1733 => "00111111",
                     1734 => "01111111",
                     1735 => "01111111",
                     1736 => "00111111",
                     1737 => "01111111",
                     1738 => "01111111",
                     1739 => "11111110",
                     1740 => "11101100",
                     1741 => "11001010",
                     1742 => "01010001",
                     1743 => "00100000",
                     1744 => "00000000",
                     1745 => "01000000",
                     1746 => "01100000",
                     1747 => "01110000",
                     1748 => "01110011",
                     1749 => "00100111",
                     1750 => "00001111",
                     1751 => "00011111",
                     1752 => "00000000",
                     1753 => "01000000",
                     1754 => "01100011",
                     1755 => "01110111",
                     1756 => "01111100",
                     1757 => "00111000",
                     1758 => "11111000",
                     1759 => "11100100",
                     1760 => "00000000",
                     1761 => "00000000",
                     1762 => "00000000",
                     1763 => "00000000",
                     1764 => "00000011",
                     1765 => "00000111",
                     1766 => "00001111",
                     1767 => "00011111",
                     1768 => "00000000",
                     1769 => "00000000",
                     1770 => "00000011",
                     1771 => "00000111",
                     1772 => "00001100",
                     1773 => "00011000",
                     1774 => "11111000",
                     1775 => "11100100",
                     1776 => "01111111",
                     1777 => "01111111",
                     1778 => "00111111",
                     1779 => "00111111",
                     1780 => "00011111",
                     1781 => "00011111",
                     1782 => "00001111",
                     1783 => "00000111",
                     1784 => "00000011",
                     1785 => "01000100",
                     1786 => "00101000",
                     1787 => "00010000",
                     1788 => "00001000",
                     1789 => "00000100",
                     1790 => "00000011",
                     1791 => "00000100",
                     1792 => "00000011",
                     1793 => "00000111",
                     1794 => "00001111",
                     1795 => "00011111",
                     1796 => "00111111",
                     1797 => "01110111",
                     1798 => "01110111",
                     1799 => "11110101",
                     1800 => "00000011",
                     1801 => "00000111",
                     1802 => "00001111",
                     1803 => "00011111",
                     1804 => "00100111",
                     1805 => "01111011",
                     1806 => "01111000",
                     1807 => "11111011",
                     1808 => "11000000",
                     1809 => "11100000",
                     1810 => "11110000",
                     1811 => "11111000",
                     1812 => "11111100",
                     1813 => "11101110",
                     1814 => "11101110",
                     1815 => "10101111",
                     1816 => "11000000",
                     1817 => "11100000",
                     1818 => "11110000",
                     1819 => "11111000",
                     1820 => "11100100",
                     1821 => "11011110",
                     1822 => "00011110",
                     1823 => "11011111",
                     1824 => "11110001",
                     1825 => "11111111",
                     1826 => "01111000",
                     1827 => "00000000",
                     1828 => "00000000",
                     1829 => "00011000",
                     1830 => "00011100",
                     1831 => "00001110",
                     1832 => "11111111",
                     1833 => "11111111",
                     1834 => "01111111",
                     1835 => "00001111",
                     1836 => "00001111",
                     1837 => "00000111",
                     1838 => "00000011",
                     1839 => "00000000",
                     1840 => "10001111",
                     1841 => "11111111",
                     1842 => "00011110",
                     1843 => "00000000",
                     1844 => "00001100",
                     1845 => "00111110",
                     1846 => "01111110",
                     1847 => "01111100",
                     1848 => "11111111",
                     1849 => "11111111",
                     1850 => "11111110",
                     1851 => "11110000",
                     1852 => "11110000",
                     1853 => "11000000",
                     1854 => "10000000",
                     1855 => "00000000",
                     1856 => "00000000",
                     1857 => "00000000",
                     1858 => "00000000",
                     1859 => "00000000",
                     1860 => "00000000",
                     1861 => "00000000",
                     1862 => "00000000",
                     1863 => "00000000",
                     1864 => "00000000",
                     1865 => "00000000",
                     1866 => "00011000",
                     1867 => "00100100",
                     1868 => "00100100",
                     1869 => "00011000",
                     1870 => "00000000",
                     1871 => "00000000",
                     1872 => "00000000",
                     1873 => "00000010",
                     1874 => "01000001",
                     1875 => "01000001",
                     1876 => "01100001",
                     1877 => "00110011",
                     1878 => "00000110",
                     1879 => "00111100",
                     1880 => "00111100",
                     1881 => "01111110",
                     1882 => "11111111",
                     1883 => "11111111",
                     1884 => "11111111",
                     1885 => "11111111",
                     1886 => "01111110",
                     1887 => "00111100",
                     1888 => "00000011",
                     1889 => "00000111",
                     1890 => "00001111",
                     1891 => "00011111",
                     1892 => "00111111",
                     1893 => "01111111",
                     1894 => "01111111",
                     1895 => "11111111",
                     1896 => "00000011",
                     1897 => "00000111",
                     1898 => "00001111",
                     1899 => "00011111",
                     1900 => "00111111",
                     1901 => "01100011",
                     1902 => "01000001",
                     1903 => "11000001",
                     1904 => "11000000",
                     1905 => "11100000",
                     1906 => "11110000",
                     1907 => "11111000",
                     1908 => "11111100",
                     1909 => "11111110",
                     1910 => "11111110",
                     1911 => "11111111",
                     1912 => "11000000",
                     1913 => "10000000",
                     1914 => "00000000",
                     1915 => "00000000",
                     1916 => "10001100",
                     1917 => "11111110",
                     1918 => "11111110",
                     1919 => "11110011",
                     1920 => "11111111",
                     1921 => "11111111",
                     1922 => "11111111",
                     1923 => "01111000",
                     1924 => "00000000",
                     1925 => "00000000",
                     1926 => "00000000",
                     1927 => "00000000",
                     1928 => "11000001",
                     1929 => "11100011",
                     1930 => "11111111",
                     1931 => "01000111",
                     1932 => "00001111",
                     1933 => "00001111",
                     1934 => "00001111",
                     1935 => "00000111",
                     1936 => "11111111",
                     1937 => "11111111",
                     1938 => "11111111",
                     1939 => "00011110",
                     1940 => "00000000",
                     1941 => "00100000",
                     1942 => "00100000",
                     1943 => "01000000",
                     1944 => "11110001",
                     1945 => "11111001",
                     1946 => "11111111",
                     1947 => "11100010",
                     1948 => "11110000",
                     1949 => "11110000",
                     1950 => "11110000",
                     1951 => "11100000",
                     1952 => "00010110",
                     1953 => "00011111",
                     1954 => "00111111",
                     1955 => "01111111",
                     1956 => "00111101",
                     1957 => "00011101",
                     1958 => "00111111",
                     1959 => "00011111",
                     1960 => "00010110",
                     1961 => "00011111",
                     1962 => "00000000",
                     1963 => "00000000",
                     1964 => "00000101",
                     1965 => "00001101",
                     1966 => "00111111",
                     1967 => "00011111",
                     1968 => "10000000",
                     1969 => "10000000",
                     1970 => "11000000",
                     1971 => "11100000",
                     1972 => "11110000",
                     1973 => "11110000",
                     1974 => "11110000",
                     1975 => "11111000",
                     1976 => "10000000",
                     1977 => "10000000",
                     1978 => "00000000",
                     1979 => "00000000",
                     1980 => "00000000",
                     1981 => "10100000",
                     1982 => "10100000",
                     1983 => "11100000",
                     1984 => "00111100",
                     1985 => "11111010",
                     1986 => "10110001",
                     1987 => "01110010",
                     1988 => "11110010",
                     1989 => "11011011",
                     1990 => "11011111",
                     1991 => "01011111",
                     1992 => "00000000",
                     1993 => "00000100",
                     1994 => "01001110",
                     1995 => "10001100",
                     1996 => "00001100",
                     1997 => "01111111",
                     1998 => "11111111",
                     1999 => "11111111",
                     2000 => "00000000",
                     2001 => "00000000",
                     2002 => "00000000",
                     2003 => "00000001",
                     2004 => "00000001",
                     2005 => "00000001",
                     2006 => "00000110",
                     2007 => "00011110",
                     2008 => "00000000",
                     2009 => "00000000",
                     2010 => "00000000",
                     2011 => "00000000",
                     2012 => "00000000",
                     2013 => "00000000",
                     2014 => "00000001",
                     2015 => "00000001",
                     2016 => "00000000",
                     2017 => "00000000",
                     2018 => "00000000",
                     2019 => "00000000",
                     2020 => "00000000",
                     2021 => "00000000",
                     2022 => "00000000",
                     2023 => "00000000",
                     2024 => "11111111",
                     2025 => "01111111",
                     2026 => "00111111",
                     2027 => "00011111",
                     2028 => "00001111",
                     2029 => "00000111",
                     2030 => "00000011",
                     2031 => "00000001",
                     2032 => "00000000",
                     2033 => "01111100",
                     2034 => "11010110",
                     2035 => "10010010",
                     2036 => "10111010",
                     2037 => "11101110",
                     2038 => "11111110",
                     2039 => "00111000",
                     2040 => "11111111",
                     2041 => "10000011",
                     2042 => "00101001",
                     2043 => "01101101",
                     2044 => "01000101",
                     2045 => "00010001",
                     2046 => "00000001",
                     2047 => "11000111",
                     2048 => "00000000",
                     2049 => "00010101",
                     2050 => "00111111",
                     2051 => "01100010",
                     2052 => "01011111",
                     2053 => "11111111",
                     2054 => "10011111",
                     2055 => "01111101",
                     2056 => "00001000",
                     2057 => "00001000",
                     2058 => "00000010",
                     2059 => "00011111",
                     2060 => "00100010",
                     2061 => "00000010",
                     2062 => "00000010",
                     2063 => "00000000",
                     2064 => "00000000",
                     2065 => "00000000",
                     2066 => "00000000",
                     2067 => "00000000",
                     2068 => "00000000",
                     2069 => "00000000",
                     2070 => "00000000",
                     2071 => "00000000",
                     2072 => "00001000",
                     2073 => "00001000",
                     2074 => "00001000",
                     2075 => "00001000",
                     2076 => "00001000",
                     2077 => "00001000",
                     2078 => "00001000",
                     2079 => "00001000",
                     2080 => "00101111",
                     2081 => "00011110",
                     2082 => "00101111",
                     2083 => "00101111",
                     2084 => "00101111",
                     2085 => "00010101",
                     2086 => "00001101",
                     2087 => "00001110",
                     2088 => "00010000",
                     2089 => "00011110",
                     2090 => "00010000",
                     2091 => "01010000",
                     2092 => "00010000",
                     2093 => "00001000",
                     2094 => "00000000",
                     2095 => "00000000",
                     2096 => "00000000",
                     2097 => "00000000",
                     2098 => "00000000",
                     2099 => "00000000",
                     2100 => "00000000",
                     2101 => "00000000",
                     2102 => "00000000",
                     2103 => "00000000",
                     2104 => "00000000",
                     2105 => "00000000",
                     2106 => "00000000",
                     2107 => "11111110",
                     2108 => "00000000",
                     2109 => "00000000",
                     2110 => "00000000",
                     2111 => "00000000",
                     2112 => "00011100",
                     2113 => "00111110",
                     2114 => "01111111",
                     2115 => "11111111",
                     2116 => "11111111",
                     2117 => "11111110",
                     2118 => "01111100",
                     2119 => "00111000",
                     2120 => "00011100",
                     2121 => "00101010",
                     2122 => "01110111",
                     2123 => "11101110",
                     2124 => "11011101",
                     2125 => "10101010",
                     2126 => "01110100",
                     2127 => "00101000",
                     2128 => "00000000",
                     2129 => "11111111",
                     2130 => "11111111",
                     2131 => "11111111",
                     2132 => "11111111",
                     2133 => "11111111",
                     2134 => "11111111",
                     2135 => "11111111",
                     2136 => "11111111",
                     2137 => "11111110",
                     2138 => "11111110",
                     2139 => "00000000",
                     2140 => "11101111",
                     2141 => "11101111",
                     2142 => "11101111",
                     2143 => "00000000",
                     2144 => "11111111",
                     2145 => "11111111",
                     2146 => "11111111",
                     2147 => "11111111",
                     2148 => "11111111",
                     2149 => "11111111",
                     2150 => "11111111",
                     2151 => "11111111",
                     2152 => "11111110",
                     2153 => "11111110",
                     2154 => "11111110",
                     2155 => "00000000",
                     2156 => "11101111",
                     2157 => "11101111",
                     2158 => "11101111",
                     2159 => "00000000",
                     2160 => "01111111",
                     2161 => "11111111",
                     2162 => "11111111",
                     2163 => "11111111",
                     2164 => "11111111",
                     2165 => "11111111",
                     2166 => "11111111",
                     2167 => "11111111",
                     2168 => "00000000",
                     2169 => "01111111",
                     2170 => "01011111",
                     2171 => "01111111",
                     2172 => "01111111",
                     2173 => "01111111",
                     2174 => "01111111",
                     2175 => "01111111",
                     2176 => "01101000",
                     2177 => "01001110",
                     2178 => "11100000",
                     2179 => "11100000",
                     2180 => "11100000",
                     2181 => "11110000",
                     2182 => "11111000",
                     2183 => "11111100",
                     2184 => "10111000",
                     2185 => "10011110",
                     2186 => "10000000",
                     2187 => "11000000",
                     2188 => "11100000",
                     2189 => "11110000",
                     2190 => "11111000",
                     2191 => "01111100",
                     2192 => "00111111",
                     2193 => "01011100",
                     2194 => "00111001",
                     2195 => "00111011",
                     2196 => "10111011",
                     2197 => "11111001",
                     2198 => "11111100",
                     2199 => "11111110",
                     2200 => "00000000",
                     2201 => "00100011",
                     2202 => "01010111",
                     2203 => "01001111",
                     2204 => "01010111",
                     2205 => "00100111",
                     2206 => "11000011",
                     2207 => "00100001",
                     2208 => "11000000",
                     2209 => "11110000",
                     2210 => "11110000",
                     2211 => "11110000",
                     2212 => "11110000",
                     2213 => "11100000",
                     2214 => "11000000",
                     2215 => "00000000",
                     2216 => "00000000",
                     2217 => "00110000",
                     2218 => "01110000",
                     2219 => "01110000",
                     2220 => "11110000",
                     2221 => "11100000",
                     2222 => "11000000",
                     2223 => "00000000",
                     2224 => "11111110",
                     2225 => "11111100",
                     2226 => "01100001",
                     2227 => "00001111",
                     2228 => "11111111",
                     2229 => "11111110",
                     2230 => "11110000",
                     2231 => "11100000",
                     2232 => "00010011",
                     2233 => "00001111",
                     2234 => "00011110",
                     2235 => "11110000",
                     2236 => "11111100",
                     2237 => "11111000",
                     2238 => "11110000",
                     2239 => "11100000",
                     2240 => "01101110",
                     2241 => "01000000",
                     2242 => "11100000",
                     2243 => "11100000",
                     2244 => "11100000",
                     2245 => "11100000",
                     2246 => "11100000",
                     2247 => "11000000",
                     2248 => "10111110",
                     2249 => "10010000",
                     2250 => "10000000",
                     2251 => "11000000",
                     2252 => "11000000",
                     2253 => "10000000",
                     2254 => "00000000",
                     2255 => "00000000",
                     2256 => "00000001",
                     2257 => "00000001",
                     2258 => "00000011",
                     2259 => "00000011",
                     2260 => "00000111",
                     2261 => "01111111",
                     2262 => "01111111",
                     2263 => "00111111",
                     2264 => "00000001",
                     2265 => "00000001",
                     2266 => "00000011",
                     2267 => "00000011",
                     2268 => "00000111",
                     2269 => "01111111",
                     2270 => "01111101",
                     2271 => "00111101",
                     2272 => "00000110",
                     2273 => "00000111",
                     2274 => "00111111",
                     2275 => "00111100",
                     2276 => "00011001",
                     2277 => "01111011",
                     2278 => "01111111",
                     2279 => "00111111",
                     2280 => "00000110",
                     2281 => "00000100",
                     2282 => "00110000",
                     2283 => "00100011",
                     2284 => "00000110",
                     2285 => "01100100",
                     2286 => "01100000",
                     2287 => "00000000",
                     2288 => "00111111",
                     2289 => "01111111",
                     2290 => "01111111",
                     2291 => "00011111",
                     2292 => "00111111",
                     2293 => "00111111",
                     2294 => "00000111",
                     2295 => "00000110",
                     2296 => "00000000",
                     2297 => "01100000",
                     2298 => "01100000",
                     2299 => "00000000",
                     2300 => "00100000",
                     2301 => "00110000",
                     2302 => "00000100",
                     2303 => "00000110",
                     2304 => "00000011",
                     2305 => "00000111",
                     2306 => "00001111",
                     2307 => "00001111",
                     2308 => "00001111",
                     2309 => "00001111",
                     2310 => "00000111",
                     2311 => "00000011",
                     2312 => "00000000",
                     2313 => "00000001",
                     2314 => "00000001",
                     2315 => "00000000",
                     2316 => "00000000",
                     2317 => "00000000",
                     2318 => "00000000",
                     2319 => "00000000",
                     2320 => "11111000",
                     2321 => "11111000",
                     2322 => "11111000",
                     2323 => "10100000",
                     2324 => "11100001",
                     2325 => "11111111",
                     2326 => "11111111",
                     2327 => "11111111",
                     2328 => "11111110",
                     2329 => "11111111",
                     2330 => "11111111",
                     2331 => "01000000",
                     2332 => "00000001",
                     2333 => "00000011",
                     2334 => "00000011",
                     2335 => "00000011",
                     2336 => "00001111",
                     2337 => "00001111",
                     2338 => "00001111",
                     2339 => "00011111",
                     2340 => "00011111",
                     2341 => "00011111",
                     2342 => "00001111",
                     2343 => "00000111",
                     2344 => "00000001",
                     2345 => "00000001",
                     2346 => "00000000",
                     2347 => "00000000",
                     2348 => "00000000",
                     2349 => "00000000",
                     2350 => "00000000",
                     2351 => "00000000",
                     2352 => "11100000",
                     2353 => "11111000",
                     2354 => "11111000",
                     2355 => "11111000",
                     2356 => "11111111",
                     2357 => "11111110",
                     2358 => "11110000",
                     2359 => "11000000",
                     2360 => "11100000",
                     2361 => "11111110",
                     2362 => "11111111",
                     2363 => "01111111",
                     2364 => "00000011",
                     2365 => "00000010",
                     2366 => "00000000",
                     2367 => "00000000",
                     2368 => "00000001",
                     2369 => "00001111",
                     2370 => "00001111",
                     2371 => "00011111",
                     2372 => "00111001",
                     2373 => "00110011",
                     2374 => "00110111",
                     2375 => "01111111",
                     2376 => "00000001",
                     2377 => "00001101",
                     2378 => "00001000",
                     2379 => "00000000",
                     2380 => "00110110",
                     2381 => "00101100",
                     2382 => "00001000",
                     2383 => "01100000",
                     2384 => "01111111",
                     2385 => "00111111",
                     2386 => "00111111",
                     2387 => "00111111",
                     2388 => "00011111",
                     2389 => "00001111",
                     2390 => "00001111",
                     2391 => "00000001",
                     2392 => "01100000",
                     2393 => "00000000",
                     2394 => "00100000",
                     2395 => "00110000",
                     2396 => "00000000",
                     2397 => "00001000",
                     2398 => "00001101",
                     2399 => "00000001",
                     2400 => "00000000",
                     2401 => "00000000",
                     2402 => "00000011",
                     2403 => "00000011",
                     2404 => "01000111",
                     2405 => "01100111",
                     2406 => "01110111",
                     2407 => "01110111",
                     2408 => "00000001",
                     2409 => "00000001",
                     2410 => "00000011",
                     2411 => "01000011",
                     2412 => "01100111",
                     2413 => "01110111",
                     2414 => "01111011",
                     2415 => "01111000",
                     2416 => "00000000",
                     2417 => "00000000",
                     2418 => "00000000",
                     2419 => "00000000",
                     2420 => "10001000",
                     2421 => "10011000",
                     2422 => "11111000",
                     2423 => "11110000",
                     2424 => "00000000",
                     2425 => "00000000",
                     2426 => "10000000",
                     2427 => "10000100",
                     2428 => "11001100",
                     2429 => "11011100",
                     2430 => "10111100",
                     2431 => "00111100",
                     2432 => "01111110",
                     2433 => "01111111",
                     2434 => "11111111",
                     2435 => "00011111",
                     2436 => "00000111",
                     2437 => "00110000",
                     2438 => "00011100",
                     2439 => "00001100",
                     2440 => "00110011",
                     2441 => "00000111",
                     2442 => "00000111",
                     2443 => "11100011",
                     2444 => "00111000",
                     2445 => "00111111",
                     2446 => "00011100",
                     2447 => "00001100",
                     2448 => "01111110",
                     2449 => "00111000",
                     2450 => "11110110",
                     2451 => "11101101",
                     2452 => "11011111",
                     2453 => "00111000",
                     2454 => "01110000",
                     2455 => "01100000",
                     2456 => "10011000",
                     2457 => "11000111",
                     2458 => "11001000",
                     2459 => "10010010",
                     2460 => "00110000",
                     2461 => "11111000",
                     2462 => "01110000",
                     2463 => "01100000",
                     2464 => "00000000",
                     2465 => "00000000",
                     2466 => "00000000",
                     2467 => "00000011",
                     2468 => "00000011",
                     2469 => "01000111",
                     2470 => "01100111",
                     2471 => "01110111",
                     2472 => "00000000",
                     2473 => "00000001",
                     2474 => "00000001",
                     2475 => "00000011",
                     2476 => "01000011",
                     2477 => "01100111",
                     2478 => "01110111",
                     2479 => "01111011",
                     2480 => "00000000",
                     2481 => "00000000",
                     2482 => "00000000",
                     2483 => "00000000",
                     2484 => "00000000",
                     2485 => "10001000",
                     2486 => "10011000",
                     2487 => "11111000",
                     2488 => "00000000",
                     2489 => "00000000",
                     2490 => "00000000",
                     2491 => "10000000",
                     2492 => "10000100",
                     2493 => "11001100",
                     2494 => "11011100",
                     2495 => "10111100",
                     2496 => "01110111",
                     2497 => "01111110",
                     2498 => "01111111",
                     2499 => "11111111",
                     2500 => "00011111",
                     2501 => "00000111",
                     2502 => "01110000",
                     2503 => "11110000",
                     2504 => "01111000",
                     2505 => "00110011",
                     2506 => "00000111",
                     2507 => "00000111",
                     2508 => "11100011",
                     2509 => "00111000",
                     2510 => "01111111",
                     2511 => "11110000",
                     2512 => "11110000",
                     2513 => "01111110",
                     2514 => "00111000",
                     2515 => "11110110",
                     2516 => "11101101",
                     2517 => "11011111",
                     2518 => "00111000",
                     2519 => "00111100",
                     2520 => "00111100",
                     2521 => "10011000",
                     2522 => "11000111",
                     2523 => "11001000",
                     2524 => "10010010",
                     2525 => "00110000",
                     2526 => "11111000",
                     2527 => "00111100",
                     2528 => "00000011",
                     2529 => "00000111",
                     2530 => "00001010",
                     2531 => "00011010",
                     2532 => "00011100",
                     2533 => "00011110",
                     2534 => "00001011",
                     2535 => "00001000",
                     2536 => "00000000",
                     2537 => "00010000",
                     2538 => "01111111",
                     2539 => "01111111",
                     2540 => "01111111",
                     2541 => "00011111",
                     2542 => "00001111",
                     2543 => "00001111",
                     2544 => "00011100",
                     2545 => "00111111",
                     2546 => "00111111",
                     2547 => "00111101",
                     2548 => "00111111",
                     2549 => "00011111",
                     2550 => "00000000",
                     2551 => "00000000",
                     2552 => "00000011",
                     2553 => "00110011",
                     2554 => "00111001",
                     2555 => "00111010",
                     2556 => "00111000",
                     2557 => "00011000",
                     2558 => "00000000",
                     2559 => "00000000",
                     2560 => "00000000",
                     2561 => "00000000",
                     2562 => "00000100",
                     2563 => "01001100",
                     2564 => "01001110",
                     2565 => "01001110",
                     2566 => "01000110",
                     2567 => "01101111",
                     2568 => "00010000",
                     2569 => "00111000",
                     2570 => "00111100",
                     2571 => "01110100",
                     2572 => "01110110",
                     2573 => "01110110",
                     2574 => "01111110",
                     2575 => "01111101",
                     2576 => "00000000",
                     2577 => "00011111",
                     2578 => "00111111",
                     2579 => "00111111",
                     2580 => "01001111",
                     2581 => "01011111",
                     2582 => "01111111",
                     2583 => "01111111",
                     2584 => "00000000",
                     2585 => "00000000",
                     2586 => "00010001",
                     2587 => "00001010",
                     2588 => "00110100",
                     2589 => "00101010",
                     2590 => "01010001",
                     2591 => "00100000",
                     2592 => "01111111",
                     2593 => "01100111",
                     2594 => "10100011",
                     2595 => "10110000",
                     2596 => "11011000",
                     2597 => "11011110",
                     2598 => "11011100",
                     2599 => "11001000",
                     2600 => "01111111",
                     2601 => "01100111",
                     2602 => "01100011",
                     2603 => "01110000",
                     2604 => "00111000",
                     2605 => "00111110",
                     2606 => "01111100",
                     2607 => "10111000",
                     2608 => "01111111",
                     2609 => "01111111",
                     2610 => "01111111",
                     2611 => "00011111",
                     2612 => "01000111",
                     2613 => "01110000",
                     2614 => "01110000",
                     2615 => "00111001",
                     2616 => "01010001",
                     2617 => "00001010",
                     2618 => "00000100",
                     2619 => "11101010",
                     2620 => "01111001",
                     2621 => "01111111",
                     2622 => "01110000",
                     2623 => "00111001",
                     2624 => "11101000",
                     2625 => "11101000",
                     2626 => "11100000",
                     2627 => "11000000",
                     2628 => "00010000",
                     2629 => "01110000",
                     2630 => "11100000",
                     2631 => "11000000",
                     2632 => "01011000",
                     2633 => "00111000",
                     2634 => "00010000",
                     2635 => "00110000",
                     2636 => "11110000",
                     2637 => "11110000",
                     2638 => "11100000",
                     2639 => "11000000",
                     2640 => "00000000",
                     2641 => "00000000",
                     2642 => "00000000",
                     2643 => "00100000",
                     2644 => "01100110",
                     2645 => "01100110",
                     2646 => "01100110",
                     2647 => "01100010",
                     2648 => "00000000",
                     2649 => "00001000",
                     2650 => "00011100",
                     2651 => "00111100",
                     2652 => "01111010",
                     2653 => "01111010",
                     2654 => "01111010",
                     2655 => "01111110",
                     2656 => "00000000",
                     2657 => "00000000",
                     2658 => "00011111",
                     2659 => "00111111",
                     2660 => "01111111",
                     2661 => "01001111",
                     2662 => "01011111",
                     2663 => "01111111",
                     2664 => "00000000",
                     2665 => "00000000",
                     2666 => "00000000",
                     2667 => "00010001",
                     2668 => "00001010",
                     2669 => "00110100",
                     2670 => "00101010",
                     2671 => "01010001",
                     2672 => "01110111",
                     2673 => "01111111",
                     2674 => "00111111",
                     2675 => "10110111",
                     2676 => "10110011",
                     2677 => "11011011",
                     2678 => "11011010",
                     2679 => "11011000",
                     2680 => "01111111",
                     2681 => "01111101",
                     2682 => "00111111",
                     2683 => "00110111",
                     2684 => "00110011",
                     2685 => "00111011",
                     2686 => "00111010",
                     2687 => "01111000",
                     2688 => "01111111",
                     2689 => "01111111",
                     2690 => "01111111",
                     2691 => "01111111",
                     2692 => "00011111",
                     2693 => "00000111",
                     2694 => "01110000",
                     2695 => "11110000",
                     2696 => "00100000",
                     2697 => "01010001",
                     2698 => "00001010",
                     2699 => "00000100",
                     2700 => "11101010",
                     2701 => "00111001",
                     2702 => "01111111",
                     2703 => "11110000",
                     2704 => "11001100",
                     2705 => "11101000",
                     2706 => "11101000",
                     2707 => "11100000",
                     2708 => "11000000",
                     2709 => "00011000",
                     2710 => "01111100",
                     2711 => "00111110",
                     2712 => "10111100",
                     2713 => "01011000",
                     2714 => "00111000",
                     2715 => "00010000",
                     2716 => "00110000",
                     2717 => "11111000",
                     2718 => "11111100",
                     2719 => "00111110",
                     2720 => "00000011",
                     2721 => "00001111",
                     2722 => "00011111",
                     2723 => "00111111",
                     2724 => "00111011",
                     2725 => "00111111",
                     2726 => "01111111",
                     2727 => "01111111",
                     2728 => "00000000",
                     2729 => "00000000",
                     2730 => "00000000",
                     2731 => "00000110",
                     2732 => "00001110",
                     2733 => "00001100",
                     2734 => "00000000",
                     2735 => "00000000",
                     2736 => "10000000",
                     2737 => "11110000",
                     2738 => "11111000",
                     2739 => "11111100",
                     2740 => "11111110",
                     2741 => "11111110",
                     2742 => "11111111",
                     2743 => "11111110",
                     2744 => "00000000",
                     2745 => "00000000",
                     2746 => "00000000",
                     2747 => "00000000",
                     2748 => "00000000",
                     2749 => "00000000",
                     2750 => "00001111",
                     2751 => "00011000",
                     2752 => "01111111",
                     2753 => "01111111",
                     2754 => "01111111",
                     2755 => "01111111",
                     2756 => "11111111",
                     2757 => "00001111",
                     2758 => "00000011",
                     2759 => "00000000",
                     2760 => "00000000",
                     2761 => "00000000",
                     2762 => "00000000",
                     2763 => "00000000",
                     2764 => "11111000",
                     2765 => "00111110",
                     2766 => "00111011",
                     2767 => "00011000",
                     2768 => "11111110",
                     2769 => "11111011",
                     2770 => "11111111",
                     2771 => "11111111",
                     2772 => "11110110",
                     2773 => "11100000",
                     2774 => "11000000",
                     2775 => "00000000",
                     2776 => "00010000",
                     2777 => "00010100",
                     2778 => "00010000",
                     2779 => "00010000",
                     2780 => "00111000",
                     2781 => "01111000",
                     2782 => "11111000",
                     2783 => "00110000",
                     2784 => "00000000",
                     2785 => "00000011",
                     2786 => "00001111",
                     2787 => "00011111",
                     2788 => "00111111",
                     2789 => "00111011",
                     2790 => "00111111",
                     2791 => "01111111",
                     2792 => "00000000",
                     2793 => "00000000",
                     2794 => "00000000",
                     2795 => "00000000",
                     2796 => "00000110",
                     2797 => "00001110",
                     2798 => "00001100",
                     2799 => "00000000",
                     2800 => "00000000",
                     2801 => "11000000",
                     2802 => "11110000",
                     2803 => "11111000",
                     2804 => "11111100",
                     2805 => "11111110",
                     2806 => "11111110",
                     2807 => "11111111",
                     2808 => "00000000",
                     2809 => "00000000",
                     2810 => "00000000",
                     2811 => "00000000",
                     2812 => "00000000",
                     2813 => "00000000",
                     2814 => "00000000",
                     2815 => "00001111",
                     2816 => "01111111",
                     2817 => "01111111",
                     2818 => "01111111",
                     2819 => "01111111",
                     2820 => "01111111",
                     2821 => "11111111",
                     2822 => "00001111",
                     2823 => "00000011",
                     2824 => "00000000",
                     2825 => "00000000",
                     2826 => "00000000",
                     2827 => "00000000",
                     2828 => "00000000",
                     2829 => "11111000",
                     2830 => "01111110",
                     2831 => "11110011",
                     2832 => "11111110",
                     2833 => "11111110",
                     2834 => "11111011",
                     2835 => "11111111",
                     2836 => "11111111",
                     2837 => "11110110",
                     2838 => "11100000",
                     2839 => "11000000",
                     2840 => "00011000",
                     2841 => "00010000",
                     2842 => "00010100",
                     2843 => "00010000",
                     2844 => "00010000",
                     2845 => "00111000",
                     2846 => "01111100",
                     2847 => "11011110",
                     2848 => "00000000",
                     2849 => "00000001",
                     2850 => "00000001",
                     2851 => "00000001",
                     2852 => "00000001",
                     2853 => "00000000",
                     2854 => "00000000",
                     2855 => "00001000",
                     2856 => "00000000",
                     2857 => "00001101",
                     2858 => "00011110",
                     2859 => "00011110",
                     2860 => "00011110",
                     2861 => "00011111",
                     2862 => "00001111",
                     2863 => "00000111",
                     2864 => "01111000",
                     2865 => "11110000",
                     2866 => "11111000",
                     2867 => "11100100",
                     2868 => "11000000",
                     2869 => "11001010",
                     2870 => "11001010",
                     2871 => "11000000",
                     2872 => "01111000",
                     2873 => "11110000",
                     2874 => "00000000",
                     2875 => "00011010",
                     2876 => "00111111",
                     2877 => "00110101",
                     2878 => "00110101",
                     2879 => "00111111",
                     2880 => "00001111",
                     2881 => "00011111",
                     2882 => "10011111",
                     2883 => "11111111",
                     2884 => "11111111",
                     2885 => "01111111",
                     2886 => "01110100",
                     2887 => "00100000",
                     2888 => "00000000",
                     2889 => "00000000",
                     2890 => "10000000",
                     2891 => "11100000",
                     2892 => "11100000",
                     2893 => "01110000",
                     2894 => "01110011",
                     2895 => "00100001",
                     2896 => "11100100",
                     2897 => "11111111",
                     2898 => "11111110",
                     2899 => "11111100",
                     2900 => "10011100",
                     2901 => "00011110",
                     2902 => "00000000",
                     2903 => "00000000",
                     2904 => "00011010",
                     2905 => "00000111",
                     2906 => "00001100",
                     2907 => "00011000",
                     2908 => "01111000",
                     2909 => "11111110",
                     2910 => "11111100",
                     2911 => "11110000",
                     2912 => "00000000",
                     2913 => "00000001",
                     2914 => "00000011",
                     2915 => "00000011",
                     2916 => "00000111",
                     2917 => "00000011",
                     2918 => "00000001",
                     2919 => "00000000",
                     2920 => "00000000",
                     2921 => "00000001",
                     2922 => "00000010",
                     2923 => "00000000",
                     2924 => "00111000",
                     2925 => "01111100",
                     2926 => "01111110",
                     2927 => "00111111",
                     2928 => "00000000",
                     2929 => "01011111",
                     2930 => "01111111",
                     2931 => "01111111",
                     2932 => "00111111",
                     2933 => "00111111",
                     2934 => "00010100",
                     2935 => "00000000",
                     2936 => "00111111",
                     2937 => "01000000",
                     2938 => "01100000",
                     2939 => "01100000",
                     2940 => "00100000",
                     2941 => "00110000",
                     2942 => "00010011",
                     2943 => "00000001",
                     2944 => "11000000",
                     2945 => "11100000",
                     2946 => "11110000",
                     2947 => "00110000",
                     2948 => "00111000",
                     2949 => "00111100",
                     2950 => "00111100",
                     2951 => "11111100",
                     2952 => "11000000",
                     2953 => "11100000",
                     2954 => "00110000",
                     2955 => "11010000",
                     2956 => "11010000",
                     2957 => "11010000",
                     2958 => "11010000",
                     2959 => "00000000",
                     2960 => "00000111",
                     2961 => "00001111",
                     2962 => "00011111",
                     2963 => "00100010",
                     2964 => "00100000",
                     2965 => "00100101",
                     2966 => "00100101",
                     2967 => "00011111",
                     2968 => "00000111",
                     2969 => "00001111",
                     2970 => "00000010",
                     2971 => "00011101",
                     2972 => "00011111",
                     2973 => "00011010",
                     2974 => "00011010",
                     2975 => "00000010",
                     2976 => "11111110",
                     2977 => "11111110",
                     2978 => "01111110",
                     2979 => "00111010",
                     2980 => "00000010",
                     2981 => "00000001",
                     2982 => "01000001",
                     2983 => "01000001",
                     2984 => "00111000",
                     2985 => "01111100",
                     2986 => "11111100",
                     2987 => "11111100",
                     2988 => "11111100",
                     2989 => "11111110",
                     2990 => "10111110",
                     2991 => "10111110",
                     2992 => "00011111",
                     2993 => "00111111",
                     2994 => "01111110",
                     2995 => "01011100",
                     2996 => "01000000",
                     2997 => "10000000",
                     2998 => "10000010",
                     2999 => "10000010",
                     3000 => "00011100",
                     3001 => "00111110",
                     3002 => "00111111",
                     3003 => "00111111",
                     3004 => "00111111",
                     3005 => "01111111",
                     3006 => "01111101",
                     3007 => "01111101",
                     3008 => "10000010",
                     3009 => "10000000",
                     3010 => "10100000",
                     3011 => "01000100",
                     3012 => "01000011",
                     3013 => "01000000",
                     3014 => "00100001",
                     3015 => "00011110",
                     3016 => "01111101",
                     3017 => "01111111",
                     3018 => "01011111",
                     3019 => "00111011",
                     3020 => "00111100",
                     3021 => "00111111",
                     3022 => "00011110",
                     3023 => "00000000",
                     3024 => "00011100",
                     3025 => "00111111",
                     3026 => "00111110",
                     3027 => "00111100",
                     3028 => "01000000",
                     3029 => "10000000",
                     3030 => "10000010",
                     3031 => "10000010",
                     3032 => "00011100",
                     3033 => "00111110",
                     3034 => "00111111",
                     3035 => "00011111",
                     3036 => "00111111",
                     3037 => "01111111",
                     3038 => "01111101",
                     3039 => "01111101",
                     3040 => "00000000",
                     3041 => "00000000",
                     3042 => "10000000",
                     3043 => "10000000",
                     3044 => "10010010",
                     3045 => "10011101",
                     3046 => "11000111",
                     3047 => "11101111",
                     3048 => "00000000",
                     3049 => "00000000",
                     3050 => "00000000",
                     3051 => "01100000",
                     3052 => "01100010",
                     3053 => "01100101",
                     3054 => "00111111",
                     3055 => "00011111",
                     3056 => "00000000",
                     3057 => "00100011",
                     3058 => "00110011",
                     3059 => "00111111",
                     3060 => "00111111",
                     3061 => "01111111",
                     3062 => "01111111",
                     3063 => "01111111",
                     3064 => "01110000",
                     3065 => "00111100",
                     3066 => "00111100",
                     3067 => "00011000",
                     3068 => "00000000",
                     3069 => "00000000",
                     3070 => "00000010",
                     3071 => "00000111",
                     3072 => "11111110",
                     3073 => "11111000",
                     3074 => "10100000",
                     3075 => "00000000",
                     3076 => "00000000",
                     3077 => "00000000",
                     3078 => "10000000",
                     3079 => "10000000",
                     3080 => "11001111",
                     3081 => "01111010",
                     3082 => "01011010",
                     3083 => "00010000",
                     3084 => "00000000",
                     3085 => "00000000",
                     3086 => "11000000",
                     3087 => "10000000",
                     3088 => "01111110",
                     3089 => "01111111",
                     3090 => "01111101",
                     3091 => "00111111",
                     3092 => "00011110",
                     3093 => "10001111",
                     3094 => "10001111",
                     3095 => "00011001",
                     3096 => "10000101",
                     3097 => "10000100",
                     3098 => "10000110",
                     3099 => "11000110",
                     3100 => "11100111",
                     3101 => "01110011",
                     3102 => "01110011",
                     3103 => "11100001",
                     3104 => "11100000",
                     3105 => "00001110",
                     3106 => "01110011",
                     3107 => "11110011",
                     3108 => "11111001",
                     3109 => "11111001",
                     3110 => "11111000",
                     3111 => "01110000",
                     3112 => "10000000",
                     3113 => "01001110",
                     3114 => "01110111",
                     3115 => "11110011",
                     3116 => "11111011",
                     3117 => "11111001",
                     3118 => "11111010",
                     3119 => "01111000",
                     3120 => "00001110",
                     3121 => "01100110",
                     3122 => "11100010",
                     3123 => "11110110",
                     3124 => "11111111",
                     3125 => "11111111",
                     3126 => "00011111",
                     3127 => "10011000",
                     3128 => "00010001",
                     3129 => "00111001",
                     3130 => "01111101",
                     3131 => "00111001",
                     3132 => "00000000",
                     3133 => "00000000",
                     3134 => "11100000",
                     3135 => "11100111",
                     3136 => "00000000",
                     3137 => "00000000",
                     3138 => "00000000",
                     3139 => "00000100",
                     3140 => "00001111",
                     3141 => "00001111",
                     3142 => "00011111",
                     3143 => "00000111",
                     3144 => "00000000",
                     3145 => "00000000",
                     3146 => "00000111",
                     3147 => "00000111",
                     3148 => "00010110",
                     3149 => "00010000",
                     3150 => "00000000",
                     3151 => "00111000",
                     3152 => "11110011",
                     3153 => "11100111",
                     3154 => "11101110",
                     3155 => "11101100",
                     3156 => "11001101",
                     3157 => "11001111",
                     3158 => "11001111",
                     3159 => "11011111",
                     3160 => "11001111",
                     3161 => "00011111",
                     3162 => "00010111",
                     3163 => "00010000",
                     3164 => "00110011",
                     3165 => "00110000",
                     3166 => "00110000",
                     3167 => "00100000",
                     3168 => "00100111",
                     3169 => "00111111",
                     3170 => "00111111",
                     3171 => "01111000",
                     3172 => "00111100",
                     3173 => "00011111",
                     3174 => "00011111",
                     3175 => "01110011",
                     3176 => "00111000",
                     3177 => "00110000",
                     3178 => "01000000",
                     3179 => "11000111",
                     3180 => "00000111",
                     3181 => "01100110",
                     3182 => "11100000",
                     3183 => "01101100",
                     3184 => "10011111",
                     3185 => "00111110",
                     3186 => "01111100",
                     3187 => "11111100",
                     3188 => "11111000",
                     3189 => "11111000",
                     3190 => "11000000",
                     3191 => "01000000",
                     3192 => "01100000",
                     3193 => "11000000",
                     3194 => "10000000",
                     3195 => "00000100",
                     3196 => "10011110",
                     3197 => "11111111",
                     3198 => "11110000",
                     3199 => "11111000",
                     3200 => "01111111",
                     3201 => "01111110",
                     3202 => "01111000",
                     3203 => "00000001",
                     3204 => "00000111",
                     3205 => "00011111",
                     3206 => "00111100",
                     3207 => "01111100",
                     3208 => "00100100",
                     3209 => "00000001",
                     3210 => "00000111",
                     3211 => "11111110",
                     3212 => "11111111",
                     3213 => "01111111",
                     3214 => "00111111",
                     3215 => "01111111",
                     3216 => "11111100",
                     3217 => "11111000",
                     3218 => "10100000",
                     3219 => "11111110",
                     3220 => "11111100",
                     3221 => "11110000",
                     3222 => "10000000",
                     3223 => "00000000",
                     3224 => "11001111",
                     3225 => "01111010",
                     3226 => "00001010",
                     3227 => "11111110",
                     3228 => "11111100",
                     3229 => "00000000",
                     3230 => "00000000",
                     3231 => "00000000",
                     3232 => "01111110",
                     3233 => "01111111",
                     3234 => "01111111",
                     3235 => "00111111",
                     3236 => "00011111",
                     3237 => "10001111",
                     3238 => "10001111",
                     3239 => "00011000",
                     3240 => "10000101",
                     3241 => "10000110",
                     3242 => "10000011",
                     3243 => "11000011",
                     3244 => "11100001",
                     3245 => "01110000",
                     3246 => "01110000",
                     3247 => "11100000",
                     3248 => "10011111",
                     3249 => "00111110",
                     3250 => "01111100",
                     3251 => "11111000",
                     3252 => "11111000",
                     3253 => "00111100",
                     3254 => "00011000",
                     3255 => "11111000",
                     3256 => "01100000",
                     3257 => "11000000",
                     3258 => "10000000",
                     3259 => "00000000",
                     3260 => "10011000",
                     3261 => "11111100",
                     3262 => "11111110",
                     3263 => "11111111",
                     3264 => "01111111",
                     3265 => "01111111",
                     3266 => "01111000",
                     3267 => "00000001",
                     3268 => "00000111",
                     3269 => "00010011",
                     3270 => "11110001",
                     3271 => "00000011",
                     3272 => "00100100",
                     3273 => "00000000",
                     3274 => "00000111",
                     3275 => "11111110",
                     3276 => "11111111",
                     3277 => "01111111",
                     3278 => "11111111",
                     3279 => "00000011",
                     3280 => "00000000",
                     3281 => "00000000",
                     3282 => "00011100",
                     3283 => "00011101",
                     3284 => "00011011",
                     3285 => "11000011",
                     3286 => "11100011",
                     3287 => "11100001",
                     3288 => "00000011",
                     3289 => "00001111",
                     3290 => "00100011",
                     3291 => "01100010",
                     3292 => "01100100",
                     3293 => "00111100",
                     3294 => "00011100",
                     3295 => "00011110",
                     3296 => "11100000",
                     3297 => "11001101",
                     3298 => "00011101",
                     3299 => "01001111",
                     3300 => "11101110",
                     3301 => "11111111",
                     3302 => "00111111",
                     3303 => "00111111",
                     3304 => "00011111",
                     3305 => "00111101",
                     3306 => "01101101",
                     3307 => "01001111",
                     3308 => "11101110",
                     3309 => "11110011",
                     3310 => "00100000",
                     3311 => "00000011",
                     3312 => "00111111",
                     3313 => "00111111",
                     3314 => "00000000",
                     3315 => "00000000",
                     3316 => "01110000",
                     3317 => "10111000",
                     3318 => "11111100",
                     3319 => "11111100",
                     3320 => "00000111",
                     3321 => "00000111",
                     3322 => "00011111",
                     3323 => "00111111",
                     3324 => "00001111",
                     3325 => "01000111",
                     3326 => "00000011",
                     3327 => "00000000",
                     3328 => "00000111",
                     3329 => "00001111",
                     3330 => "00011111",
                     3331 => "00111111",
                     3332 => "00111110",
                     3333 => "01111100",
                     3334 => "01111000",
                     3335 => "01111000",
                     3336 => "00000000",
                     3337 => "00000000",
                     3338 => "00000011",
                     3339 => "00000111",
                     3340 => "00001111",
                     3341 => "00001111",
                     3342 => "00011111",
                     3343 => "00011111",
                     3344 => "00111111",
                     3345 => "01011100",
                     3346 => "00111001",
                     3347 => "00111011",
                     3348 => "10111111",
                     3349 => "11111111",
                     3350 => "11111110",
                     3351 => "11111110",
                     3352 => "00000000",
                     3353 => "00100011",
                     3354 => "01010111",
                     3355 => "01001111",
                     3356 => "01010111",
                     3357 => "00101111",
                     3358 => "11011111",
                     3359 => "00100001",
                     3360 => "11000000",
                     3361 => "11000000",
                     3362 => "10000000",
                     3363 => "10000000",
                     3364 => "10000000",
                     3365 => "10000000",
                     3366 => "00000000",
                     3367 => "00000000",
                     3368 => "00000000",
                     3369 => "00000000",
                     3370 => "00000000",
                     3371 => "00000000",
                     3372 => "10000000",
                     3373 => "10000000",
                     3374 => "00000000",
                     3375 => "00000000",
                     3376 => "11111110",
                     3377 => "11111100",
                     3378 => "01100001",
                     3379 => "00001111",
                     3380 => "01111111",
                     3381 => "00111111",
                     3382 => "00011111",
                     3383 => "00011110",
                     3384 => "00100011",
                     3385 => "00001111",
                     3386 => "00011110",
                     3387 => "11110000",
                     3388 => "00011100",
                     3389 => "00111111",
                     3390 => "00011111",
                     3391 => "00011110",
                     3392 => "11110000",
                     3393 => "01111000",
                     3394 => "11100100",
                     3395 => "11001000",
                     3396 => "11001100",
                     3397 => "10111110",
                     3398 => "10111110",
                     3399 => "00111110",
                     3400 => "00000000",
                     3401 => "10000000",
                     3402 => "00011000",
                     3403 => "00110000",
                     3404 => "00110100",
                     3405 => "11111110",
                     3406 => "11111110",
                     3407 => "11111110",
                     3408 => "00000000",
                     3409 => "00000001",
                     3410 => "00000000",
                     3411 => "00000111",
                     3412 => "00000111",
                     3413 => "00000111",
                     3414 => "00000111",
                     3415 => "00011111",
                     3416 => "00000000",
                     3417 => "00000000",
                     3418 => "00000001",
                     3419 => "00000100",
                     3420 => "00000110",
                     3421 => "00000110",
                     3422 => "00000111",
                     3423 => "00000111",
                     3424 => "00000000",
                     3425 => "00000000",
                     3426 => "00001111",
                     3427 => "00111111",
                     3428 => "00111111",
                     3429 => "00001111",
                     3430 => "00000000",
                     3431 => "00000000",
                     3432 => "00001111",
                     3433 => "00111111",
                     3434 => "01111111",
                     3435 => "11111000",
                     3436 => "11111000",
                     3437 => "01111111",
                     3438 => "00111111",
                     3439 => "00001111",
                     3440 => "01111000",
                     3441 => "01111100",
                     3442 => "01111110",
                     3443 => "01111111",
                     3444 => "00111111",
                     3445 => "00111111",
                     3446 => "00011011",
                     3447 => "00001001",
                     3448 => "00011111",
                     3449 => "00011111",
                     3450 => "00011111",
                     3451 => "00001011",
                     3452 => "00000001",
                     3453 => "00000001",
                     3454 => "00000000",
                     3455 => "00000000",
                     3456 => "00001100",
                     3457 => "00000000",
                     3458 => "00000000",
                     3459 => "00000000",
                     3460 => "00000111",
                     3461 => "01111111",
                     3462 => "01111100",
                     3463 => "00000000",
                     3464 => "00000011",
                     3465 => "00011111",
                     3466 => "00111111",
                     3467 => "00111111",
                     3468 => "01111000",
                     3469 => "00000000",
                     3470 => "00000011",
                     3471 => "11111111",
                     3472 => "00000001",
                     3473 => "11100001",
                     3474 => "01110001",
                     3475 => "01111001",
                     3476 => "00111101",
                     3477 => "00111101",
                     3478 => "00011111",
                     3479 => "00000011",
                     3480 => "00000000",
                     3481 => "00000000",
                     3482 => "00000000",
                     3483 => "00000000",
                     3484 => "00000000",
                     3485 => "00000000",
                     3486 => "00000000",
                     3487 => "00000000",
                     3488 => "00111111",
                     3489 => "00111111",
                     3490 => "00011111",
                     3491 => "00011011",
                     3492 => "00110110",
                     3493 => "00110000",
                     3494 => "01111111",
                     3495 => "00111111",
                     3496 => "00100011",
                     3497 => "00100111",
                     3498 => "00011111",
                     3499 => "00000111",
                     3500 => "00001111",
                     3501 => "00011111",
                     3502 => "01111111",
                     3503 => "00111111",
                     3504 => "11111000",
                     3505 => "11111000",
                     3506 => "11111000",
                     3507 => "10111000",
                     3508 => "00011000",
                     3509 => "11011000",
                     3510 => "11011000",
                     3511 => "10111000",
                     3512 => "11100000",
                     3513 => "10000000",
                     3514 => "10000000",
                     3515 => "01000000",
                     3516 => "11100000",
                     3517 => "11100000",
                     3518 => "11100000",
                     3519 => "11000000",
                     3520 => "00000001",
                     3521 => "00000010",
                     3522 => "00000100",
                     3523 => "00000100",
                     3524 => "00001000",
                     3525 => "00001000",
                     3526 => "00010000",
                     3527 => "00010000",
                     3528 => "00000011",
                     3529 => "00000111",
                     3530 => "00001111",
                     3531 => "00011111",
                     3532 => "00111111",
                     3533 => "01111111",
                     3534 => "11111111",
                     3535 => "00011111",
                     3536 => "00000000",
                     3537 => "00001111",
                     3538 => "00010011",
                     3539 => "00001101",
                     3540 => "00001101",
                     3541 => "00010011",
                     3542 => "00001100",
                     3543 => "00100000",
                     3544 => "00011111",
                     3545 => "00010000",
                     3546 => "00001100",
                     3547 => "00010010",
                     3548 => "00010010",
                     3549 => "00101100",
                     3550 => "00111111",
                     3551 => "00111111",
                     3552 => "00000000",
                     3553 => "00100100",
                     3554 => "00000000",
                     3555 => "00100100",
                     3556 => "00000000",
                     3557 => "00000100",
                     3558 => "00000000",
                     3559 => "00000000",
                     3560 => "00110111",
                     3561 => "00110110",
                     3562 => "00110110",
                     3563 => "00110110",
                     3564 => "00010110",
                     3565 => "00010110",
                     3566 => "00010010",
                     3567 => "00000010",
                     3568 => "00001111",
                     3569 => "01000001",
                     3570 => "00000000",
                     3571 => "10001000",
                     3572 => "00000000",
                     3573 => "01000100",
                     3574 => "00000000",
                     3575 => "00000000",
                     3576 => "00010000",
                     3577 => "01111110",
                     3578 => "11111111",
                     3579 => "11111111",
                     3580 => "11110110",
                     3581 => "01110110",
                     3582 => "00111010",
                     3583 => "00011010",
                     3584 => "00111000",
                     3585 => "01111100",
                     3586 => "11111110",
                     3587 => "11111110",
                     3588 => "00111011",
                     3589 => "00000011",
                     3590 => "00000011",
                     3591 => "00000011",
                     3592 => "00000000",
                     3593 => "00000000",
                     3594 => "00111000",
                     3595 => "00000100",
                     3596 => "00000000",
                     3597 => "00000000",
                     3598 => "00000000",
                     3599 => "00000000",
                     3600 => "00000011",
                     3601 => "00110011",
                     3602 => "01111011",
                     3603 => "01111111",
                     3604 => "11111111",
                     3605 => "11111011",
                     3606 => "00000011",
                     3607 => "00000011",
                     3608 => "00000000",
                     3609 => "00000000",
                     3610 => "00000000",
                     3611 => "00111000",
                     3612 => "01000000",
                     3613 => "00000000",
                     3614 => "00000000",
                     3615 => "00000000",
                     3616 => "11011100",
                     3617 => "11000000",
                     3618 => "11100000",
                     3619 => "11100000",
                     3620 => "11100000",
                     3621 => "11100000",
                     3622 => "11100000",
                     3623 => "11000000",
                     3624 => "11111100",
                     3625 => "10100000",
                     3626 => "10000000",
                     3627 => "10000000",
                     3628 => "00000000",
                     3629 => "00000000",
                     3630 => "00000000",
                     3631 => "00000000",
                     3632 => "00111111",
                     3633 => "01011111",
                     3634 => "00111111",
                     3635 => "00111111",
                     3636 => "10111011",
                     3637 => "11111000",
                     3638 => "11111110",
                     3639 => "11111110",
                     3640 => "00000111",
                     3641 => "00100111",
                     3642 => "01010111",
                     3643 => "01001111",
                     3644 => "01010111",
                     3645 => "00100111",
                     3646 => "11000001",
                     3647 => "00100001",
                     3648 => "00011111",
                     3649 => "00001111",
                     3650 => "00001111",
                     3651 => "00011111",
                     3652 => "00011111",
                     3653 => "00011110",
                     3654 => "00111000",
                     3655 => "00110000",
                     3656 => "00011101",
                     3657 => "00001111",
                     3658 => "00001111",
                     3659 => "00011111",
                     3660 => "00011111",
                     3661 => "00011110",
                     3662 => "00111000",
                     3663 => "00110000",
                     3664 => "00000000",
                     3665 => "00100000",
                     3666 => "01100000",
                     3667 => "01100000",
                     3668 => "01110000",
                     3669 => "11110000",
                     3670 => "11111000",
                     3671 => "11111000",
                     3672 => "00000000",
                     3673 => "00000000",
                     3674 => "00111000",
                     3675 => "00010000",
                     3676 => "01001100",
                     3677 => "00011000",
                     3678 => "10000110",
                     3679 => "00100100",
                     3680 => "11111000",
                     3681 => "11111100",
                     3682 => "11111100",
                     3683 => "01111110",
                     3684 => "01111110",
                     3685 => "00111110",
                     3686 => "00011111",
                     3687 => "00000111",
                     3688 => "00000000",
                     3689 => "01000010",
                     3690 => "00001010",
                     3691 => "01000000",
                     3692 => "00010000",
                     3693 => "00000010",
                     3694 => "00001000",
                     3695 => "00000010",
                     3696 => "00000000",
                     3697 => "11000000",
                     3698 => "01110000",
                     3699 => "10111000",
                     3700 => "11110100",
                     3701 => "11110010",
                     3702 => "11110101",
                     3703 => "01111011",
                     3704 => "00000000",
                     3705 => "00000000",
                     3706 => "10000000",
                     3707 => "01000000",
                     3708 => "00001000",
                     3709 => "00001100",
                     3710 => "00001010",
                     3711 => "10000100",
                     3712 => "00000000",
                     3713 => "11011111",
                     3714 => "00010000",
                     3715 => "11111111",
                     3716 => "11011111",
                     3717 => "11111111",
                     3718 => "11111111",
                     3719 => "11111001",
                     3720 => "00000000",
                     3721 => "00000000",
                     3722 => "11001111",
                     3723 => "00100000",
                     3724 => "00100000",
                     3725 => "00100000",
                     3726 => "00100110",
                     3727 => "00101110",
                     3728 => "00011111",
                     3729 => "00011111",
                     3730 => "00111110",
                     3731 => "11111100",
                     3732 => "11111000",
                     3733 => "11110000",
                     3734 => "11000000",
                     3735 => "00000000",
                     3736 => "11100000",
                     3737 => "11100000",
                     3738 => "11000000",
                     3739 => "00000000",
                     3740 => "00000000",
                     3741 => "00000000",
                     3742 => "00000000",
                     3743 => "00000000",
                     3744 => "11111000",
                     3745 => "11111100",
                     3746 => "11111110",
                     3747 => "11111111",
                     3748 => "11111111",
                     3749 => "11011111",
                     3750 => "11011111",
                     3751 => "00000000",
                     3752 => "00101111",
                     3753 => "00100011",
                     3754 => "00100001",
                     3755 => "00100000",
                     3756 => "00100000",
                     3757 => "00000000",
                     3758 => "00000000",
                     3759 => "00000000",
                     3760 => "11000001",
                     3761 => "11110001",
                     3762 => "01111001",
                     3763 => "01111101",
                     3764 => "00111101",
                     3765 => "00111111",
                     3766 => "00011111",
                     3767 => "00000011",
                     3768 => "11000001",
                     3769 => "10110001",
                     3770 => "01011001",
                     3771 => "01101101",
                     3772 => "00110101",
                     3773 => "00111011",
                     3774 => "00011111",
                     3775 => "00000011",
                     3776 => "00000010",
                     3777 => "00000110",
                     3778 => "00001110",
                     3779 => "00001110",
                     3780 => "00011110",
                     3781 => "00011110",
                     3782 => "00111110",
                     3783 => "00111110",
                     3784 => "00000000",
                     3785 => "00000010",
                     3786 => "00000000",
                     3787 => "00001000",
                     3788 => "00000010",
                     3789 => "00000000",
                     3790 => "00101000",
                     3791 => "00000000",
                     3792 => "00111110",
                     3793 => "00111110",
                     3794 => "00111110",
                     3795 => "00111110",
                     3796 => "00011110",
                     3797 => "00011110",
                     3798 => "00001110",
                     3799 => "00000010",
                     3800 => "00000100",
                     3801 => "00010000",
                     3802 => "00000010",
                     3803 => "00010000",
                     3804 => "00000100",
                     3805 => "00000000",
                     3806 => "00001010",
                     3807 => "00000000",
                     3808 => "11000001",
                     3809 => "11110001",
                     3810 => "01111001",
                     3811 => "01111101",
                     3812 => "00111101",
                     3813 => "00111111",
                     3814 => "00011111",
                     3815 => "00000011",
                     3816 => "11000001",
                     3817 => "10110001",
                     3818 => "01011001",
                     3819 => "01101101",
                     3820 => "00110101",
                     3821 => "00111011",
                     3822 => "00011111",
                     3823 => "00000011",
                     3824 => "01111100",
                     3825 => "00000000",
                     3826 => "00000000",
                     3827 => "11111111",
                     3828 => "11000011",
                     3829 => "01111111",
                     3830 => "00011111",
                     3831 => "00000011",
                     3832 => "00000000",
                     3833 => "00001111",
                     3834 => "00011111",
                     3835 => "11111111",
                     3836 => "11111100",
                     3837 => "01100011",
                     3838 => "00011111",
                     3839 => "00000011",
                     3840 => "11111111",
                     3841 => "11111111",
                     3842 => "01111100",
                     3843 => "00000000",
                     3844 => "00000000",
                     3845 => "01111100",
                     3846 => "11111111",
                     3847 => "11111111",
                     3848 => "00000000",
                     3849 => "00000000",
                     3850 => "11111110",
                     3851 => "11000110",
                     3852 => "11000110",
                     3853 => "11111110",
                     3854 => "00000000",
                     3855 => "00000000",
                     3856 => "11111111",
                     3857 => "11111111",
                     3858 => "00000000",
                     3859 => "00000100",
                     3860 => "00001100",
                     3861 => "00011000",
                     3862 => "00110000",
                     3863 => "00000000",
                     3864 => "00000000",
                     3865 => "00000000",
                     3866 => "00000110",
                     3867 => "00000110",
                     3868 => "00001100",
                     3869 => "00011000",
                     3870 => "01110000",
                     3871 => "01100000",
                     3872 => "11111111",
                     3873 => "11111111",
                     3874 => "00000000",
                     3875 => "00000100",
                     3876 => "00000100",
                     3877 => "00000100",
                     3878 => "00001000",
                     3879 => "00001000",
                     3880 => "00000000",
                     3881 => "00000000",
                     3882 => "00000110",
                     3883 => "00000110",
                     3884 => "00000100",
                     3885 => "00000100",
                     3886 => "00001000",
                     3887 => "00001000",
                     3888 => "00001000",
                     3889 => "00010000",
                     3890 => "00010000",
                     3891 => "00000000",
                     3892 => "00000000",
                     3893 => "00010000",
                     3894 => "00010000",
                     3895 => "00001000",
                     3896 => "00001000",
                     3897 => "00010000",
                     3898 => "00110000",
                     3899 => "00110000",
                     3900 => "00110000",
                     3901 => "00110000",
                     3902 => "00010000",
                     3903 => "00001000",
                     3904 => "01111111",
                     3905 => "00111111",
                     3906 => "00111111",
                     3907 => "00111110",
                     3908 => "00011111",
                     3909 => "00001111",
                     3910 => "00000011",
                     3911 => "00000000",
                     3912 => "00000000",
                     3913 => "00000000",
                     3914 => "00000001",
                     3915 => "00000011",
                     3916 => "00000001",
                     3917 => "00000000",
                     3918 => "00000000",
                     3919 => "00000000",
                     3920 => "00000011",
                     3921 => "00001111",
                     3922 => "11111111",
                     3923 => "01111111",
                     3924 => "01111111",
                     3925 => "01111111",
                     3926 => "01111111",
                     3927 => "01111111",
                     3928 => "00000011",
                     3929 => "00001110",
                     3930 => "11111000",
                     3931 => "00000000",
                     3932 => "00000000",
                     3933 => "00000000",
                     3934 => "00000000",
                     3935 => "00000000",
                     3936 => "00000000",
                     3937 => "00000000",
                     3938 => "00000000",
                     3939 => "00000000",
                     3940 => "00000000",
                     3941 => "00000000",
                     3942 => "00000000",
                     3943 => "00000000",
                     3944 => "00100010",
                     3945 => "01100101",
                     3946 => "00100101",
                     3947 => "00100101",
                     3948 => "00100101",
                     3949 => "00100101",
                     3950 => "01110111",
                     3951 => "01110010",
                     3952 => "00000000",
                     3953 => "00000000",
                     3954 => "00000000",
                     3955 => "00000000",
                     3956 => "00000000",
                     3957 => "00000000",
                     3958 => "00000000",
                     3959 => "00000000",
                     3960 => "01100010",
                     3961 => "10010101",
                     3962 => "00010101",
                     3963 => "00100101",
                     3964 => "01000101",
                     3965 => "10000101",
                     3966 => "11110111",
                     3967 => "11110010",
                     3968 => "00000000",
                     3969 => "00000000",
                     3970 => "00000000",
                     3971 => "00000000",
                     3972 => "00000000",
                     3973 => "00000000",
                     3974 => "00000000",
                     3975 => "00000000",
                     3976 => "10100010",
                     3977 => "10100101",
                     3978 => "10100101",
                     3979 => "10100101",
                     3980 => "11110101",
                     3981 => "11110101",
                     3982 => "00100111",
                     3983 => "00100010",
                     3984 => "00000000",
                     3985 => "00000000",
                     3986 => "00000000",
                     3987 => "00000000",
                     3988 => "00000000",
                     3989 => "00000000",
                     3990 => "00000000",
                     3991 => "00000000",
                     3992 => "11110010",
                     3993 => "10000101",
                     3994 => "10000101",
                     3995 => "11100101",
                     3996 => "00010101",
                     3997 => "00010101",
                     3998 => "11110111",
                     3999 => "11100010",
                     4000 => "00000000",
                     4001 => "00000000",
                     4002 => "00000000",
                     4003 => "00000000",
                     4004 => "00000000",
                     4005 => "00000000",
                     4006 => "00000000",
                     4007 => "00000000",
                     4008 => "01100010",
                     4009 => "10010101",
                     4010 => "01010101",
                     4011 => "01100101",
                     4012 => "10110101",
                     4013 => "10010101",
                     4014 => "10010111",
                     4015 => "01100010",
                     4016 => "00000000",
                     4017 => "00000000",
                     4018 => "00000000",
                     4019 => "00000000",
                     4020 => "00000000",
                     4021 => "00000000",
                     4022 => "00000000",
                     4023 => "00000000",
                     4024 => "00100000",
                     4025 => "01010000",
                     4026 => "01010000",
                     4027 => "01010000",
                     4028 => "01010000",
                     4029 => "01010000",
                     4030 => "01110000",
                     4031 => "00100000",
                     4032 => "00000000",
                     4033 => "00000000",
                     4034 => "00000000",
                     4035 => "00000000",
                     4036 => "00000000",
                     4037 => "00000000",
                     4038 => "00000000",
                     4039 => "00000000",
                     4040 => "00000000",
                     4041 => "00000000",
                     4042 => "00000000",
                     4043 => "00000000",
                     4044 => "00000000",
                     4045 => "00000000",
                     4046 => "00000000",
                     4047 => "00000000",
                     4048 => "00000000",
                     4049 => "00000000",
                     4050 => "00000000",
                     4051 => "00000000",
                     4052 => "00000000",
                     4053 => "00000000",
                     4054 => "00000000",
                     4055 => "00000000",
                     4056 => "01100110",
                     4057 => "11100110",
                     4058 => "01100110",
                     4059 => "01100110",
                     4060 => "01100110",
                     4061 => "01100111",
                     4062 => "11110011",
                     4063 => "00000000",
                     4064 => "00000000",
                     4065 => "00000000",
                     4066 => "00000000",
                     4067 => "00000000",
                     4068 => "00000000",
                     4069 => "00000000",
                     4070 => "00000000",
                     4071 => "00000000",
                     4072 => "01011110",
                     4073 => "01011001",
                     4074 => "01011001",
                     4075 => "01011001",
                     4076 => "01011110",
                     4077 => "11011000",
                     4078 => "10011000",
                     4079 => "00000000",
                     4080 => "00000000",
                     4081 => "00000000",
                     4082 => "00000000",
                     4083 => "00000000",
                     4084 => "00000000",
                     4085 => "01111100",
                     4086 => "00111000",
                     4087 => "00000000",
                     4088 => "00000000",
                     4089 => "00000000",
                     4090 => "00000000",
                     4091 => "00000000",
                     4092 => "00000000",
                     4093 => "00000100",
                     4094 => "00001000",
                     4095 => "00000000",
                     4096 => "00111000",
                     4097 => "01001100",
                     4098 => "11000110",
                     4099 => "11000110",
                     4100 => "11000110",
                     4101 => "01100100",
                     4102 => "00111000",
                     4103 => "00000000",
                     4104 => "00000000",
                     4105 => "00000000",
                     4106 => "00000000",
                     4107 => "00000000",
                     4108 => "00000000",
                     4109 => "00000000",
                     4110 => "00000000",
                     4111 => "00000000",
                     4112 => "00011000",
                     4113 => "00111000",
                     4114 => "00011000",
                     4115 => "00011000",
                     4116 => "00011000",
                     4117 => "00011000",
                     4118 => "01111110",
                     4119 => "00000000",
                     4120 => "00000000",
                     4121 => "00000000",
                     4122 => "00000000",
                     4123 => "00000000",
                     4124 => "00000000",
                     4125 => "00000000",
                     4126 => "00000000",
                     4127 => "00000000",
                     4128 => "01111100",
                     4129 => "11000110",
                     4130 => "00001110",
                     4131 => "00111100",
                     4132 => "01111000",
                     4133 => "11100000",
                     4134 => "11111110",
                     4135 => "00000000",
                     4136 => "00000000",
                     4137 => "00000000",
                     4138 => "00000000",
                     4139 => "00000000",
                     4140 => "00000000",
                     4141 => "00000000",
                     4142 => "00000000",
                     4143 => "00000000",
                     4144 => "01111110",
                     4145 => "00001100",
                     4146 => "00011000",
                     4147 => "00111100",
                     4148 => "00000110",
                     4149 => "11000110",
                     4150 => "01111100",
                     4151 => "00000000",
                     4152 => "00000000",
                     4153 => "00000000",
                     4154 => "00000000",
                     4155 => "00000000",
                     4156 => "00000000",
                     4157 => "00000000",
                     4158 => "00000000",
                     4159 => "00000000",
                     4160 => "00011100",
                     4161 => "00111100",
                     4162 => "01101100",
                     4163 => "11001100",
                     4164 => "11111110",
                     4165 => "00001100",
                     4166 => "00001100",
                     4167 => "00000000",
                     4168 => "00000000",
                     4169 => "00000000",
                     4170 => "00000000",
                     4171 => "00000000",
                     4172 => "00000000",
                     4173 => "00000000",
                     4174 => "00000000",
                     4175 => "00000000",
                     4176 => "11111100",
                     4177 => "11000000",
                     4178 => "11111100",
                     4179 => "00000110",
                     4180 => "00000110",
                     4181 => "11000110",
                     4182 => "01111100",
                     4183 => "00000000",
                     4184 => "00000000",
                     4185 => "00000000",
                     4186 => "00000000",
                     4187 => "00000000",
                     4188 => "00000000",
                     4189 => "00000000",
                     4190 => "00000000",
                     4191 => "00000000",
                     4192 => "00111100",
                     4193 => "01100000",
                     4194 => "11000000",
                     4195 => "11111100",
                     4196 => "11000110",
                     4197 => "11000110",
                     4198 => "01111100",
                     4199 => "00000000",
                     4200 => "00000000",
                     4201 => "00000000",
                     4202 => "00000000",
                     4203 => "00000000",
                     4204 => "00000000",
                     4205 => "00000000",
                     4206 => "00000000",
                     4207 => "00000000",
                     4208 => "11111110",
                     4209 => "11000110",
                     4210 => "00001100",
                     4211 => "00011000",
                     4212 => "00110000",
                     4213 => "00110000",
                     4214 => "00110000",
                     4215 => "00000000",
                     4216 => "00000000",
                     4217 => "00000000",
                     4218 => "00000000",
                     4219 => "00000000",
                     4220 => "00000000",
                     4221 => "00000000",
                     4222 => "00000000",
                     4223 => "00000000",
                     4224 => "01111100",
                     4225 => "11000110",
                     4226 => "11000110",
                     4227 => "01111100",
                     4228 => "11000110",
                     4229 => "11000110",
                     4230 => "01111100",
                     4231 => "00000000",
                     4232 => "00000000",
                     4233 => "00000000",
                     4234 => "00000000",
                     4235 => "00000000",
                     4236 => "00000000",
                     4237 => "00000000",
                     4238 => "00000000",
                     4239 => "00000000",
                     4240 => "01111100",
                     4241 => "11000110",
                     4242 => "11000110",
                     4243 => "01111110",
                     4244 => "00000110",
                     4245 => "00001100",
                     4246 => "01111000",
                     4247 => "00000000",
                     4248 => "00000000",
                     4249 => "00000000",
                     4250 => "00000000",
                     4251 => "00000000",
                     4252 => "00000000",
                     4253 => "00000000",
                     4254 => "00000000",
                     4255 => "00000000",
                     4256 => "00111000",
                     4257 => "01101100",
                     4258 => "11000110",
                     4259 => "11000110",
                     4260 => "11111110",
                     4261 => "11000110",
                     4262 => "11000110",
                     4263 => "00000000",
                     4264 => "00000000",
                     4265 => "00000000",
                     4266 => "00000000",
                     4267 => "00000000",
                     4268 => "00000000",
                     4269 => "00000000",
                     4270 => "00000000",
                     4271 => "00000000",
                     4272 => "11111100",
                     4273 => "11000110",
                     4274 => "11000110",
                     4275 => "11111100",
                     4276 => "11000110",
                     4277 => "11000110",
                     4278 => "11111100",
                     4279 => "00000000",
                     4280 => "00000000",
                     4281 => "00000000",
                     4282 => "00000000",
                     4283 => "00000000",
                     4284 => "00000000",
                     4285 => "00000000",
                     4286 => "00000000",
                     4287 => "00000000",
                     4288 => "00111100",
                     4289 => "01100110",
                     4290 => "11000000",
                     4291 => "11000000",
                     4292 => "11000000",
                     4293 => "01100110",
                     4294 => "00111100",
                     4295 => "00000000",
                     4296 => "00000000",
                     4297 => "00000000",
                     4298 => "00000000",
                     4299 => "00000000",
                     4300 => "00000000",
                     4301 => "00000000",
                     4302 => "00000000",
                     4303 => "00000000",
                     4304 => "11111000",
                     4305 => "11001100",
                     4306 => "11000110",
                     4307 => "11000110",
                     4308 => "11000110",
                     4309 => "11001100",
                     4310 => "11111000",
                     4311 => "00000000",
                     4312 => "00000000",
                     4313 => "00000000",
                     4314 => "00000000",
                     4315 => "00000000",
                     4316 => "00000000",
                     4317 => "00000000",
                     4318 => "00000000",
                     4319 => "00000000",
                     4320 => "11111110",
                     4321 => "11000000",
                     4322 => "11000000",
                     4323 => "11111100",
                     4324 => "11000000",
                     4325 => "11000000",
                     4326 => "11111110",
                     4327 => "00000000",
                     4328 => "00000000",
                     4329 => "00000000",
                     4330 => "00000000",
                     4331 => "00000000",
                     4332 => "00000000",
                     4333 => "00000000",
                     4334 => "00000000",
                     4335 => "00000000",
                     4336 => "11111110",
                     4337 => "11000000",
                     4338 => "11000000",
                     4339 => "11111100",
                     4340 => "11000000",
                     4341 => "11000000",
                     4342 => "11000000",
                     4343 => "00000000",
                     4344 => "00000000",
                     4345 => "00000000",
                     4346 => "00000000",
                     4347 => "00000000",
                     4348 => "00000000",
                     4349 => "00000000",
                     4350 => "00000000",
                     4351 => "00000000",
                     4352 => "00111110",
                     4353 => "01100000",
                     4354 => "11000000",
                     4355 => "11001110",
                     4356 => "11000110",
                     4357 => "01100110",
                     4358 => "00111110",
                     4359 => "00000000",
                     4360 => "00000000",
                     4361 => "00000000",
                     4362 => "00000000",
                     4363 => "00000000",
                     4364 => "00000000",
                     4365 => "00000000",
                     4366 => "00000000",
                     4367 => "00000000",
                     4368 => "11000110",
                     4369 => "11000110",
                     4370 => "11000110",
                     4371 => "11111110",
                     4372 => "11000110",
                     4373 => "11000110",
                     4374 => "11000110",
                     4375 => "00000000",
                     4376 => "00000000",
                     4377 => "00000000",
                     4378 => "00000000",
                     4379 => "00000000",
                     4380 => "00000000",
                     4381 => "00000000",
                     4382 => "00000000",
                     4383 => "00000000",
                     4384 => "01111110",
                     4385 => "00011000",
                     4386 => "00011000",
                     4387 => "00011000",
                     4388 => "00011000",
                     4389 => "00011000",
                     4390 => "01111110",
                     4391 => "00000000",
                     4392 => "00000000",
                     4393 => "00000000",
                     4394 => "00000000",
                     4395 => "00000000",
                     4396 => "00000000",
                     4397 => "00000000",
                     4398 => "00000000",
                     4399 => "00000000",
                     4400 => "00011110",
                     4401 => "00000110",
                     4402 => "00000110",
                     4403 => "00000110",
                     4404 => "11000110",
                     4405 => "11000110",
                     4406 => "01111100",
                     4407 => "00000000",
                     4408 => "00000000",
                     4409 => "00000000",
                     4410 => "00000000",
                     4411 => "00000000",
                     4412 => "00000000",
                     4413 => "00000000",
                     4414 => "00000000",
                     4415 => "00000000",
                     4416 => "11000110",
                     4417 => "11001100",
                     4418 => "11011000",
                     4419 => "11110000",
                     4420 => "11111000",
                     4421 => "11011100",
                     4422 => "11001110",
                     4423 => "00000000",
                     4424 => "00000000",
                     4425 => "00000000",
                     4426 => "00000000",
                     4427 => "00000000",
                     4428 => "00000000",
                     4429 => "00000000",
                     4430 => "00000000",
                     4431 => "00000000",
                     4432 => "01100000",
                     4433 => "01100000",
                     4434 => "01100000",
                     4435 => "01100000",
                     4436 => "01100000",
                     4437 => "01100000",
                     4438 => "01111110",
                     4439 => "00000000",
                     4440 => "00000000",
                     4441 => "00000000",
                     4442 => "00000000",
                     4443 => "00000000",
                     4444 => "00000000",
                     4445 => "00000000",
                     4446 => "00000000",
                     4447 => "00000000",
                     4448 => "11000110",
                     4449 => "11101110",
                     4450 => "11111110",
                     4451 => "11111110",
                     4452 => "11010110",
                     4453 => "11000110",
                     4454 => "11000110",
                     4455 => "00000000",
                     4456 => "00000000",
                     4457 => "00000000",
                     4458 => "00000000",
                     4459 => "00000000",
                     4460 => "00000000",
                     4461 => "00000000",
                     4462 => "00000000",
                     4463 => "00000000",
                     4464 => "11000110",
                     4465 => "11100110",
                     4466 => "11110110",
                     4467 => "11111110",
                     4468 => "11011110",
                     4469 => "11001110",
                     4470 => "11000110",
                     4471 => "00000000",
                     4472 => "00000000",
                     4473 => "00000000",
                     4474 => "00000000",
                     4475 => "00000000",
                     4476 => "00000000",
                     4477 => "00000000",
                     4478 => "00000000",
                     4479 => "00000000",
                     4480 => "01111100",
                     4481 => "11000110",
                     4482 => "11000110",
                     4483 => "11000110",
                     4484 => "11000110",
                     4485 => "11000110",
                     4486 => "01111100",
                     4487 => "00000000",
                     4488 => "00000000",
                     4489 => "00000000",
                     4490 => "00000000",
                     4491 => "00000000",
                     4492 => "00000000",
                     4493 => "00000000",
                     4494 => "00000000",
                     4495 => "00000000",
                     4496 => "11111100",
                     4497 => "11000110",
                     4498 => "11000110",
                     4499 => "11000110",
                     4500 => "11111100",
                     4501 => "11000000",
                     4502 => "11000000",
                     4503 => "00000000",
                     4504 => "00000000",
                     4505 => "00000000",
                     4506 => "00000000",
                     4507 => "00000000",
                     4508 => "00000000",
                     4509 => "00000000",
                     4510 => "00000000",
                     4511 => "00000000",
                     4512 => "01111100",
                     4513 => "11000110",
                     4514 => "11000110",
                     4515 => "11000110",
                     4516 => "11011110",
                     4517 => "11001100",
                     4518 => "01111010",
                     4519 => "00000000",
                     4520 => "00000000",
                     4521 => "00000000",
                     4522 => "00000000",
                     4523 => "00000000",
                     4524 => "00000000",
                     4525 => "00000000",
                     4526 => "00000000",
                     4527 => "00000000",
                     4528 => "11111100",
                     4529 => "11000110",
                     4530 => "11000110",
                     4531 => "11001110",
                     4532 => "11111000",
                     4533 => "11011100",
                     4534 => "11001110",
                     4535 => "00000000",
                     4536 => "00000000",
                     4537 => "00000000",
                     4538 => "00000000",
                     4539 => "00000000",
                     4540 => "00000000",
                     4541 => "00000000",
                     4542 => "00000000",
                     4543 => "00000000",
                     4544 => "01111000",
                     4545 => "11001100",
                     4546 => "11000000",
                     4547 => "01111100",
                     4548 => "00000110",
                     4549 => "11000110",
                     4550 => "01111100",
                     4551 => "00000000",
                     4552 => "00000000",
                     4553 => "00000000",
                     4554 => "00000000",
                     4555 => "00000000",
                     4556 => "00000000",
                     4557 => "00000000",
                     4558 => "00000000",
                     4559 => "00000000",
                     4560 => "01111110",
                     4561 => "00011000",
                     4562 => "00011000",
                     4563 => "00011000",
                     4564 => "00011000",
                     4565 => "00011000",
                     4566 => "00011000",
                     4567 => "00000000",
                     4568 => "00000000",
                     4569 => "00000000",
                     4570 => "00000000",
                     4571 => "00000000",
                     4572 => "00000000",
                     4573 => "00000000",
                     4574 => "00000000",
                     4575 => "00000000",
                     4576 => "11000110",
                     4577 => "11000110",
                     4578 => "11000110",
                     4579 => "11000110",
                     4580 => "11000110",
                     4581 => "11000110",
                     4582 => "01111100",
                     4583 => "00000000",
                     4584 => "00000000",
                     4585 => "00000000",
                     4586 => "00000000",
                     4587 => "00000000",
                     4588 => "00000000",
                     4589 => "00000000",
                     4590 => "00000000",
                     4591 => "00000000",
                     4592 => "11000110",
                     4593 => "11000110",
                     4594 => "11000110",
                     4595 => "11101110",
                     4596 => "01111100",
                     4597 => "00111000",
                     4598 => "00010000",
                     4599 => "00000000",
                     4600 => "00000000",
                     4601 => "00000000",
                     4602 => "00000000",
                     4603 => "00000000",
                     4604 => "00000000",
                     4605 => "00000000",
                     4606 => "00000000",
                     4607 => "00000000",
                     4608 => "11000110",
                     4609 => "11000110",
                     4610 => "11010110",
                     4611 => "11111110",
                     4612 => "11111110",
                     4613 => "11101110",
                     4614 => "11000110",
                     4615 => "00000000",
                     4616 => "00000000",
                     4617 => "00000000",
                     4618 => "00000000",
                     4619 => "00000000",
                     4620 => "00000000",
                     4621 => "00000000",
                     4622 => "00000000",
                     4623 => "00000000",
                     4624 => "11000110",
                     4625 => "11101110",
                     4626 => "01111100",
                     4627 => "00111000",
                     4628 => "01111100",
                     4629 => "11101110",
                     4630 => "11000110",
                     4631 => "00000000",
                     4632 => "00000000",
                     4633 => "00000000",
                     4634 => "00000000",
                     4635 => "00000000",
                     4636 => "00000000",
                     4637 => "00000000",
                     4638 => "00000000",
                     4639 => "00000000",
                     4640 => "01100110",
                     4641 => "01100110",
                     4642 => "01100110",
                     4643 => "00111100",
                     4644 => "00011000",
                     4645 => "00011000",
                     4646 => "00011000",
                     4647 => "00000000",
                     4648 => "00000000",
                     4649 => "00000000",
                     4650 => "00000000",
                     4651 => "00000000",
                     4652 => "00000000",
                     4653 => "00000000",
                     4654 => "00000000",
                     4655 => "00000000",
                     4656 => "11111110",
                     4657 => "00001110",
                     4658 => "00011100",
                     4659 => "00111000",
                     4660 => "01110000",
                     4661 => "11100000",
                     4662 => "11111110",
                     4663 => "00000000",
                     4664 => "00000000",
                     4665 => "00000000",
                     4666 => "00000000",
                     4667 => "00000000",
                     4668 => "00000000",
                     4669 => "00000000",
                     4670 => "00000000",
                     4671 => "00000000",
                     4672 => "00000000",
                     4673 => "00000000",
                     4674 => "00000000",
                     4675 => "00000000",
                     4676 => "00000000",
                     4677 => "00000000",
                     4678 => "00000000",
                     4679 => "00000000",
                     4680 => "00000000",
                     4681 => "00000000",
                     4682 => "00000000",
                     4683 => "00000000",
                     4684 => "00000000",
                     4685 => "00000000",
                     4686 => "00000000",
                     4687 => "00000000",
                     4688 => "11111111",
                     4689 => "11111111",
                     4690 => "11111111",
                     4691 => "11111111",
                     4692 => "11111111",
                     4693 => "11111111",
                     4694 => "11111111",
                     4695 => "11111111",
                     4696 => "00000000",
                     4697 => "00000000",
                     4698 => "00000000",
                     4699 => "00000000",
                     4700 => "00000000",
                     4701 => "00000000",
                     4702 => "00000000",
                     4703 => "00000000",
                     4704 => "00000000",
                     4705 => "00000000",
                     4706 => "00000000",
                     4707 => "00000000",
                     4708 => "00000000",
                     4709 => "00000000",
                     4710 => "00000000",
                     4711 => "00000000",
                     4712 => "11111111",
                     4713 => "11111111",
                     4714 => "11111111",
                     4715 => "11111111",
                     4716 => "11111111",
                     4717 => "11111111",
                     4718 => "11111111",
                     4719 => "11111111",
                     4720 => "11111111",
                     4721 => "11111111",
                     4722 => "11111111",
                     4723 => "11111111",
                     4724 => "11111111",
                     4725 => "11111111",
                     4726 => "11111111",
                     4727 => "11111111",
                     4728 => "11111111",
                     4729 => "11111111",
                     4730 => "11111111",
                     4731 => "11111111",
                     4732 => "11111111",
                     4733 => "11111111",
                     4734 => "11111111",
                     4735 => "11111111",
                     4736 => "00000000",
                     4737 => "00000000",
                     4738 => "00000000",
                     4739 => "01111110",
                     4740 => "01111110",
                     4741 => "00000000",
                     4742 => "00000000",
                     4743 => "00000000",
                     4744 => "00000000",
                     4745 => "00000000",
                     4746 => "00000000",
                     4747 => "00000000",
                     4748 => "00000000",
                     4749 => "00000000",
                     4750 => "00000000",
                     4751 => "00000000",
                     4752 => "00000000",
                     4753 => "00000000",
                     4754 => "01000100",
                     4755 => "00101000",
                     4756 => "00010000",
                     4757 => "00101000",
                     4758 => "01000100",
                     4759 => "00000000",
                     4760 => "00000000",
                     4761 => "00000000",
                     4762 => "00000000",
                     4763 => "00000000",
                     4764 => "00000000",
                     4765 => "00000000",
                     4766 => "00000000",
                     4767 => "00000000",
                     4768 => "11111111",
                     4769 => "11111111",
                     4770 => "11111111",
                     4771 => "11111111",
                     4772 => "11111111",
                     4773 => "11111111",
                     4774 => "11111111",
                     4775 => "11111111",
                     4776 => "01111111",
                     4777 => "01111111",
                     4778 => "01111111",
                     4779 => "01111111",
                     4780 => "01111111",
                     4781 => "01111111",
                     4782 => "01111111",
                     4783 => "01111111",
                     4784 => "00011000",
                     4785 => "00111100",
                     4786 => "00111100",
                     4787 => "00111100",
                     4788 => "00011000",
                     4789 => "00011000",
                     4790 => "00000000",
                     4791 => "00011000",
                     4792 => "00000000",
                     4793 => "00000000",
                     4794 => "00000000",
                     4795 => "00000000",
                     4796 => "00000000",
                     4797 => "00000000",
                     4798 => "00000000",
                     4799 => "00000000",
                     4800 => "11111111",
                     4801 => "01111111",
                     4802 => "01111111",
                     4803 => "01111111",
                     4804 => "01111111",
                     4805 => "11111111",
                     4806 => "11100011",
                     4807 => "11000001",
                     4808 => "11111111",
                     4809 => "10000000",
                     4810 => "10000000",
                     4811 => "10000000",
                     4812 => "10000000",
                     4813 => "00000000",
                     4814 => "00011100",
                     4815 => "00111110",
                     4816 => "10000000",
                     4817 => "10000000",
                     4818 => "10000000",
                     4819 => "11000001",
                     4820 => "11100011",
                     4821 => "11111111",
                     4822 => "11111111",
                     4823 => "11111111",
                     4824 => "01111111",
                     4825 => "01111111",
                     4826 => "01111111",
                     4827 => "00111110",
                     4828 => "00011100",
                     4829 => "00000000",
                     4830 => "00000000",
                     4831 => "11111111",
                     4832 => "00111000",
                     4833 => "01111100",
                     4834 => "01111100",
                     4835 => "01111100",
                     4836 => "01111100",
                     4837 => "01111100",
                     4838 => "00111000",
                     4839 => "00000000",
                     4840 => "00001000",
                     4841 => "00000100",
                     4842 => "00000100",
                     4843 => "00000100",
                     4844 => "00000100",
                     4845 => "00000100",
                     4846 => "00001000",
                     4847 => "00000000",
                     4848 => "00000011",
                     4849 => "00000110",
                     4850 => "00001100",
                     4851 => "00001100",
                     4852 => "00001000",
                     4853 => "00001000",
                     4854 => "00000100",
                     4855 => "00000011",
                     4856 => "00000011",
                     4857 => "00000101",
                     4858 => "00001011",
                     4859 => "00001011",
                     4860 => "00001111",
                     4861 => "00001111",
                     4862 => "00000111",
                     4863 => "00000011",
                     4864 => "00000001",
                     4865 => "00000010",
                     4866 => "00000100",
                     4867 => "00001000",
                     4868 => "00010000",
                     4869 => "00100000",
                     4870 => "01000000",
                     4871 => "10000000",
                     4872 => "00000001",
                     4873 => "00000011",
                     4874 => "00000111",
                     4875 => "00001111",
                     4876 => "00011111",
                     4877 => "00111111",
                     4878 => "01111111",
                     4879 => "11111111",
                     4880 => "00000000",
                     4881 => "00000000",
                     4882 => "00000000",
                     4883 => "00000000",
                     4884 => "00000000",
                     4885 => "00000111",
                     4886 => "00111000",
                     4887 => "11000000",
                     4888 => "00000000",
                     4889 => "00000000",
                     4890 => "00000000",
                     4891 => "00000000",
                     4892 => "00000000",
                     4893 => "00000111",
                     4894 => "00111111",
                     4895 => "11111111",
                     4896 => "00000000",
                     4897 => "00000000",
                     4898 => "00000000",
                     4899 => "00000000",
                     4900 => "00000000",
                     4901 => "11100000",
                     4902 => "00011100",
                     4903 => "00000011",
                     4904 => "00000000",
                     4905 => "00000000",
                     4906 => "00000000",
                     4907 => "00000000",
                     4908 => "00000000",
                     4909 => "11100000",
                     4910 => "11111100",
                     4911 => "11111111",
                     4912 => "10000000",
                     4913 => "01000000",
                     4914 => "00100000",
                     4915 => "00010000",
                     4916 => "00001000",
                     4917 => "00000100",
                     4918 => "00000010",
                     4919 => "00000001",
                     4920 => "10000000",
                     4921 => "11000000",
                     4922 => "11100000",
                     4923 => "11110000",
                     4924 => "11111000",
                     4925 => "11111100",
                     4926 => "11111110",
                     4927 => "11111111",
                     4928 => "00000100",
                     4929 => "00001110",
                     4930 => "00001110",
                     4931 => "00001110",
                     4932 => "01101110",
                     4933 => "01100100",
                     4934 => "01100000",
                     4935 => "01100000",
                     4936 => "11111111",
                     4937 => "11111111",
                     4938 => "11111111",
                     4939 => "11111111",
                     4940 => "11111111",
                     4941 => "11111111",
                     4942 => "11111111",
                     4943 => "11111111",
                     4944 => "00000111",
                     4945 => "00001111",
                     4946 => "00011111",
                     4947 => "00011111",
                     4948 => "01111111",
                     4949 => "11111111",
                     4950 => "11111111",
                     4951 => "01111111",
                     4952 => "00000111",
                     4953 => "00001000",
                     4954 => "00010000",
                     4955 => "00000000",
                     4956 => "01100000",
                     4957 => "10000000",
                     4958 => "10000000",
                     4959 => "01000000",
                     4960 => "00000011",
                     4961 => "00000111",
                     4962 => "00011111",
                     4963 => "00111111",
                     4964 => "00111111",
                     4965 => "00111111",
                     4966 => "01111001",
                     4967 => "11110111",
                     4968 => "00000011",
                     4969 => "00000100",
                     4970 => "00011000",
                     4971 => "00100000",
                     4972 => "00100000",
                     4973 => "00100000",
                     4974 => "01000110",
                     4975 => "10001000",
                     4976 => "11000000",
                     4977 => "11100000",
                     4978 => "11110000",
                     4979 => "11110100",
                     4980 => "11111110",
                     4981 => "10111111",
                     4982 => "11011111",
                     4983 => "11111111",
                     4984 => "11000000",
                     4985 => "00100000",
                     4986 => "00010000",
                     4987 => "00010100",
                     4988 => "00001010",
                     4989 => "01000001",
                     4990 => "00100001",
                     4991 => "00000001",
                     4992 => "10010000",
                     4993 => "10111000",
                     4994 => "11111000",
                     4995 => "11111010",
                     4996 => "11111111",
                     4997 => "11111111",
                     4998 => "11111111",
                     4999 => "11111110",
                     5000 => "10010000",
                     5001 => "10101000",
                     5002 => "01001000",
                     5003 => "00001010",
                     5004 => "00000101",
                     5005 => "00000001",
                     5006 => "00000001",
                     5007 => "00000010",
                     5008 => "00111011",
                     5009 => "00011101",
                     5010 => "00001110",
                     5011 => "00001111",
                     5012 => "00000111",
                     5013 => "00000000",
                     5014 => "00000000",
                     5015 => "00000000",
                     5016 => "00100100",
                     5017 => "00010010",
                     5018 => "00001001",
                     5019 => "00001000",
                     5020 => "00000111",
                     5021 => "00000000",
                     5022 => "00000000",
                     5023 => "00000000",
                     5024 => "11111111",
                     5025 => "10111111",
                     5026 => "00011100",
                     5027 => "11000000",
                     5028 => "11110011",
                     5029 => "11111111",
                     5030 => "01111110",
                     5031 => "00011100",
                     5032 => "00000000",
                     5033 => "01000000",
                     5034 => "11100011",
                     5035 => "00111111",
                     5036 => "00001100",
                     5037 => "10000001",
                     5038 => "01100010",
                     5039 => "00011100",
                     5040 => "10111111",
                     5041 => "01111111",
                     5042 => "00111101",
                     5043 => "10000011",
                     5044 => "11000111",
                     5045 => "11111111",
                     5046 => "11111111",
                     5047 => "00111100",
                     5048 => "01000000",
                     5049 => "10000000",
                     5050 => "11000010",
                     5051 => "01111100",
                     5052 => "00111000",
                     5053 => "00000000",
                     5054 => "11000011",
                     5055 => "00111100",
                     5056 => "11111100",
                     5057 => "11111110",
                     5058 => "11111111",
                     5059 => "11111110",
                     5060 => "11111110",
                     5061 => "11111000",
                     5062 => "01100000",
                     5063 => "00000000",
                     5064 => "00000100",
                     5065 => "00000010",
                     5066 => "00000001",
                     5067 => "00000000",
                     5068 => "00000110",
                     5069 => "10011000",
                     5070 => "01100000",
                     5071 => "00000000",
                     5072 => "11000000",
                     5073 => "00100000",
                     5074 => "00010000",
                     5075 => "00010000",
                     5076 => "00010000",
                     5077 => "00010000",
                     5078 => "00100000",
                     5079 => "11000000",
                     5080 => "11000000",
                     5081 => "11100000",
                     5082 => "11110000",
                     5083 => "11110000",
                     5084 => "11110000",
                     5085 => "11110000",
                     5086 => "11100000",
                     5087 => "11000000",
                     5088 => "00000000",
                     5089 => "00000000",
                     5090 => "00000000",
                     5091 => "00000000",
                     5092 => "00111111",
                     5093 => "01111111",
                     5094 => "11100000",
                     5095 => "11000000",
                     5096 => "00000000",
                     5097 => "00000000",
                     5098 => "00000000",
                     5099 => "00000000",
                     5100 => "00000000",
                     5101 => "00000000",
                     5102 => "00011100",
                     5103 => "00111110",
                     5104 => "10001000",
                     5105 => "10011100",
                     5106 => "10001000",
                     5107 => "10000000",
                     5108 => "10000000",
                     5109 => "10000000",
                     5110 => "10000000",
                     5111 => "10000000",
                     5112 => "01111111",
                     5113 => "01111111",
                     5114 => "01111111",
                     5115 => "00111110",
                     5116 => "00011100",
                     5117 => "00000000",
                     5118 => "00000000",
                     5119 => "00000000",
                     5120 => "11111110",
                     5121 => "11111110",
                     5122 => "11111110",
                     5123 => "11111110",
                     5124 => "11111110",
                     5125 => "11111110",
                     5126 => "11111110",
                     5127 => "11111110",
                     5128 => "11111111",
                     5129 => "11111111",
                     5130 => "11111111",
                     5131 => "11111111",
                     5132 => "11111111",
                     5133 => "11111111",
                     5134 => "11111111",
                     5135 => "11111111",
                     5136 => "00001000",
                     5137 => "00010100",
                     5138 => "00100100",
                     5139 => "11000100",
                     5140 => "00000011",
                     5141 => "01000000",
                     5142 => "10100001",
                     5143 => "00100110",
                     5144 => "00000000",
                     5145 => "00001000",
                     5146 => "00011000",
                     5147 => "00111000",
                     5148 => "11111100",
                     5149 => "10111111",
                     5150 => "01011110",
                     5151 => "11011001",
                     5152 => "11111111",
                     5153 => "11111111",
                     5154 => "11111111",
                     5155 => "11111111",
                     5156 => "01111111",
                     5157 => "01111111",
                     5158 => "01111111",
                     5159 => "01111111",
                     5160 => "10000001",
                     5161 => "10000001",
                     5162 => "10000001",
                     5163 => "10000001",
                     5164 => "10000001",
                     5165 => "10000001",
                     5166 => "10000001",
                     5167 => "10000001",
                     5168 => "11111111",
                     5169 => "11111111",
                     5170 => "11111111",
                     5171 => "11111111",
                     5172 => "11111111",
                     5173 => "11111111",
                     5174 => "11111111",
                     5175 => "11111111",
                     5176 => "00000001",
                     5177 => "00000001",
                     5178 => "00000001",
                     5179 => "00000001",
                     5180 => "00000001",
                     5181 => "00000001",
                     5182 => "00000001",
                     5183 => "00000001",
                     5184 => "01111111",
                     5185 => "10000000",
                     5186 => "10000000",
                     5187 => "10011000",
                     5188 => "10011100",
                     5189 => "10001100",
                     5190 => "10000000",
                     5191 => "10000000",
                     5192 => "00000000",
                     5193 => "01111111",
                     5194 => "01111111",
                     5195 => "01100111",
                     5196 => "01100111",
                     5197 => "01111111",
                     5198 => "01111111",
                     5199 => "01111111",
                     5200 => "11111111",
                     5201 => "00000001",
                     5202 => "00000001",
                     5203 => "11111111",
                     5204 => "00010000",
                     5205 => "00010000",
                     5206 => "00010000",
                     5207 => "11111111",
                     5208 => "00000000",
                     5209 => "11111111",
                     5210 => "11111111",
                     5211 => "11111111",
                     5212 => "11111111",
                     5213 => "11111111",
                     5214 => "11111111",
                     5215 => "11111111",
                     5216 => "10000000",
                     5217 => "10000000",
                     5218 => "10000000",
                     5219 => "10000000",
                     5220 => "10000000",
                     5221 => "10000000",
                     5222 => "10000000",
                     5223 => "10000000",
                     5224 => "01111111",
                     5225 => "01111111",
                     5226 => "01111111",
                     5227 => "01111111",
                     5228 => "01111111",
                     5229 => "01111111",
                     5230 => "01111111",
                     5231 => "01111111",
                     5232 => "00000001",
                     5233 => "00000001",
                     5234 => "00000001",
                     5235 => "11111111",
                     5236 => "00010000",
                     5237 => "00010000",
                     5238 => "00010000",
                     5239 => "11111111",
                     5240 => "11111111",
                     5241 => "11111111",
                     5242 => "11111111",
                     5243 => "11111111",
                     5244 => "11111111",
                     5245 => "11111111",
                     5246 => "11111111",
                     5247 => "11111111",
                     5248 => "11111111",
                     5249 => "00000000",
                     5250 => "00000000",
                     5251 => "00000000",
                     5252 => "00000000",
                     5253 => "00000000",
                     5254 => "00000000",
                     5255 => "00000000",
                     5256 => "00000000",
                     5257 => "11111111",
                     5258 => "11111111",
                     5259 => "11111111",
                     5260 => "11111111",
                     5261 => "11111111",
                     5262 => "11111111",
                     5263 => "11111111",
                     5264 => "11111110",
                     5265 => "00000001",
                     5266 => "00000001",
                     5267 => "00011001",
                     5268 => "00011101",
                     5269 => "00001101",
                     5270 => "00000001",
                     5271 => "00000001",
                     5272 => "00000000",
                     5273 => "11111111",
                     5274 => "11111111",
                     5275 => "11100111",
                     5276 => "11100111",
                     5277 => "11111111",
                     5278 => "11111111",
                     5279 => "11111111",
                     5280 => "00000001",
                     5281 => "00000001",
                     5282 => "00000001",
                     5283 => "00000001",
                     5284 => "00000001",
                     5285 => "00000001",
                     5286 => "00000001",
                     5287 => "00000001",
                     5288 => "11111111",
                     5289 => "11111111",
                     5290 => "11111111",
                     5291 => "11111111",
                     5292 => "11111111",
                     5293 => "11111111",
                     5294 => "11111111",
                     5295 => "11111111",
                     5296 => "00111111",
                     5297 => "01111111",
                     5298 => "01111111",
                     5299 => "11111111",
                     5300 => "11111111",
                     5301 => "11111111",
                     5302 => "11111111",
                     5303 => "11111111",
                     5304 => "00111111",
                     5305 => "01100000",
                     5306 => "01000000",
                     5307 => "11000000",
                     5308 => "10000000",
                     5309 => "10000000",
                     5310 => "10000000",
                     5311 => "10000000",
                     5312 => "11111111",
                     5313 => "11111111",
                     5314 => "11111111",
                     5315 => "11111111",
                     5316 => "11111111",
                     5317 => "11111111",
                     5318 => "01111110",
                     5319 => "00111100",
                     5320 => "10000000",
                     5321 => "10000000",
                     5322 => "10000000",
                     5323 => "10000000",
                     5324 => "10000000",
                     5325 => "10000001",
                     5326 => "01000010",
                     5327 => "00111100",
                     5328 => "11111111",
                     5329 => "11111111",
                     5330 => "11111111",
                     5331 => "11111111",
                     5332 => "11111111",
                     5333 => "11111111",
                     5334 => "11111111",
                     5335 => "11111111",
                     5336 => "11111111",
                     5337 => "00000000",
                     5338 => "00000000",
                     5339 => "00000000",
                     5340 => "00000000",
                     5341 => "00000000",
                     5342 => "00000000",
                     5343 => "00000000",
                     5344 => "11111111",
                     5345 => "11111111",
                     5346 => "11111111",
                     5347 => "11111111",
                     5348 => "11111111",
                     5349 => "11111111",
                     5350 => "11111110",
                     5351 => "01111100",
                     5352 => "00000000",
                     5353 => "00000000",
                     5354 => "00000000",
                     5355 => "00000000",
                     5356 => "00000000",
                     5357 => "00000001",
                     5358 => "10000010",
                     5359 => "01111100",
                     5360 => "11111111",
                     5361 => "11111111",
                     5362 => "11111111",
                     5363 => "11111111",
                     5364 => "11111111",
                     5365 => "11111111",
                     5366 => "11111110",
                     5367 => "01111100",
                     5368 => "00000000",
                     5369 => "00000000",
                     5370 => "00000000",
                     5371 => "00000000",
                     5372 => "00000000",
                     5373 => "00000001",
                     5374 => "10000011",
                     5375 => "11111111",
                     5376 => "11111000",
                     5377 => "11111100",
                     5378 => "11111110",
                     5379 => "11111110",
                     5380 => "11111111",
                     5381 => "11111111",
                     5382 => "11111111",
                     5383 => "11111111",
                     5384 => "11111000",
                     5385 => "00000100",
                     5386 => "00000010",
                     5387 => "00000010",
                     5388 => "00000001",
                     5389 => "00000001",
                     5390 => "00000001",
                     5391 => "00000001",
                     5392 => "11111111",
                     5393 => "11111111",
                     5394 => "11111111",
                     5395 => "11111111",
                     5396 => "11111111",
                     5397 => "11111111",
                     5398 => "01111110",
                     5399 => "00111100",
                     5400 => "00000001",
                     5401 => "00000001",
                     5402 => "00000001",
                     5403 => "00000001",
                     5404 => "00000001",
                     5405 => "10000001",
                     5406 => "01000010",
                     5407 => "00111100",
                     5408 => "00000000",
                     5409 => "00001000",
                     5410 => "00001000",
                     5411 => "00001000",
                     5412 => "00010000",
                     5413 => "00010000",
                     5414 => "00010000",
                     5415 => "00000000",
                     5416 => "11111111",
                     5417 => "11111111",
                     5418 => "11111111",
                     5419 => "11111111",
                     5420 => "11111111",
                     5421 => "11111111",
                     5422 => "11111111",
                     5423 => "11111111",
                     5424 => "00000000",
                     5425 => "01111111",
                     5426 => "01111111",
                     5427 => "01111000",
                     5428 => "01110011",
                     5429 => "01110011",
                     5430 => "01110011",
                     5431 => "01111111",
                     5432 => "01111111",
                     5433 => "10000000",
                     5434 => "10100000",
                     5435 => "10000111",
                     5436 => "10001111",
                     5437 => "10001110",
                     5438 => "10001110",
                     5439 => "10000110",
                     5440 => "00000000",
                     5441 => "11111111",
                     5442 => "11111111",
                     5443 => "00111111",
                     5444 => "10011111",
                     5445 => "10011111",
                     5446 => "10011111",
                     5447 => "00011111",
                     5448 => "11111110",
                     5449 => "00000001",
                     5450 => "00000101",
                     5451 => "11000001",
                     5452 => "11100001",
                     5453 => "01110001",
                     5454 => "01110001",
                     5455 => "11110001",
                     5456 => "01111110",
                     5457 => "01111110",
                     5458 => "01111111",
                     5459 => "01111110",
                     5460 => "01111110",
                     5461 => "01111111",
                     5462 => "01111111",
                     5463 => "11111111",
                     5464 => "10000001",
                     5465 => "10000001",
                     5466 => "10000000",
                     5467 => "10000001",
                     5468 => "10000001",
                     5469 => "10100000",
                     5470 => "10000000",
                     5471 => "11111111",
                     5472 => "01111111",
                     5473 => "01111111",
                     5474 => "11111111",
                     5475 => "01111111",
                     5476 => "01111111",
                     5477 => "11111111",
                     5478 => "11111111",
                     5479 => "11111111",
                     5480 => "11110001",
                     5481 => "11000001",
                     5482 => "11000001",
                     5483 => "10000001",
                     5484 => "11000001",
                     5485 => "11000101",
                     5486 => "00000001",
                     5487 => "11111111",
                     5488 => "01111111",
                     5489 => "10000000",
                     5490 => "10100000",
                     5491 => "10000000",
                     5492 => "10000000",
                     5493 => "10000000",
                     5494 => "10000000",
                     5495 => "10000000",
                     5496 => "01111111",
                     5497 => "11111111",
                     5498 => "11111111",
                     5499 => "11111111",
                     5500 => "11111111",
                     5501 => "11111111",
                     5502 => "11111111",
                     5503 => "11111111",
                     5504 => "11111110",
                     5505 => "00000001",
                     5506 => "00000101",
                     5507 => "00000001",
                     5508 => "00000001",
                     5509 => "00000001",
                     5510 => "00000001",
                     5511 => "00000001",
                     5512 => "11111110",
                     5513 => "11111111",
                     5514 => "11111111",
                     5515 => "11111111",
                     5516 => "11111111",
                     5517 => "11111111",
                     5518 => "11111111",
                     5519 => "11111111",
                     5520 => "10000000",
                     5521 => "10000000",
                     5522 => "10000000",
                     5523 => "10000000",
                     5524 => "10000000",
                     5525 => "10100000",
                     5526 => "10000000",
                     5527 => "01111111",
                     5528 => "11111111",
                     5529 => "11111111",
                     5530 => "11111111",
                     5531 => "11111111",
                     5532 => "11111111",
                     5533 => "11111111",
                     5534 => "11111111",
                     5535 => "01111111",
                     5536 => "00000001",
                     5537 => "00000001",
                     5538 => "00000001",
                     5539 => "00000001",
                     5540 => "00000001",
                     5541 => "00000101",
                     5542 => "00000001",
                     5543 => "11111110",
                     5544 => "11111111",
                     5545 => "11111111",
                     5546 => "11111111",
                     5547 => "11111111",
                     5548 => "11111111",
                     5549 => "11111111",
                     5550 => "11111111",
                     5551 => "11111110",
                     5552 => "00000000",
                     5553 => "00000000",
                     5554 => "00000000",
                     5555 => "00000000",
                     5556 => "11111100",
                     5557 => "11111110",
                     5558 => "00000111",
                     5559 => "00000011",
                     5560 => "00000000",
                     5561 => "00000000",
                     5562 => "00000000",
                     5563 => "00000000",
                     5564 => "00000000",
                     5565 => "00000000",
                     5566 => "00111000",
                     5567 => "01111100",
                     5568 => "00010001",
                     5569 => "00111001",
                     5570 => "00010001",
                     5571 => "00000001",
                     5572 => "00000001",
                     5573 => "00000001",
                     5574 => "00000001",
                     5575 => "00000001",
                     5576 => "11111110",
                     5577 => "11111110",
                     5578 => "11111110",
                     5579 => "01111100",
                     5580 => "00111000",
                     5581 => "00000000",
                     5582 => "00000000",
                     5583 => "00000000",
                     5584 => "11101111",
                     5585 => "00101000",
                     5586 => "00101000",
                     5587 => "00101000",
                     5588 => "00101000",
                     5589 => "00101000",
                     5590 => "11101111",
                     5591 => "00000000",
                     5592 => "00100000",
                     5593 => "11100111",
                     5594 => "11100111",
                     5595 => "11100111",
                     5596 => "11100111",
                     5597 => "11100111",
                     5598 => "11101111",
                     5599 => "00000000",
                     5600 => "11111110",
                     5601 => "10000010",
                     5602 => "10000010",
                     5603 => "10000010",
                     5604 => "10000010",
                     5605 => "10000010",
                     5606 => "11111110",
                     5607 => "00000000",
                     5608 => "00000010",
                     5609 => "01111110",
                     5610 => "01111110",
                     5611 => "01111110",
                     5612 => "01111110",
                     5613 => "01111110",
                     5614 => "11111110",
                     5615 => "00000000",
                     5616 => "10000000",
                     5617 => "10000000",
                     5618 => "10000000",
                     5619 => "10011000",
                     5620 => "10011100",
                     5621 => "10001100",
                     5622 => "10000000",
                     5623 => "01111111",
                     5624 => "01111111",
                     5625 => "01111111",
                     5626 => "01111111",
                     5627 => "01100111",
                     5628 => "01100111",
                     5629 => "01111111",
                     5630 => "01111111",
                     5631 => "01111111",
                     5632 => "11111111",
                     5633 => "11111111",
                     5634 => "10000011",
                     5635 => "11110011",
                     5636 => "11110011",
                     5637 => "11110011",
                     5638 => "11110011",
                     5639 => "11110011",
                     5640 => "11111111",
                     5641 => "10000000",
                     5642 => "11111100",
                     5643 => "10001100",
                     5644 => "10001100",
                     5645 => "10001100",
                     5646 => "10001100",
                     5647 => "10001100",
                     5648 => "11111111",
                     5649 => "11111111",
                     5650 => "11110000",
                     5651 => "11110110",
                     5652 => "11110110",
                     5653 => "11110110",
                     5654 => "11110110",
                     5655 => "11110110",
                     5656 => "11111111",
                     5657 => "00000000",
                     5658 => "00001111",
                     5659 => "00001001",
                     5660 => "00001001",
                     5661 => "00001001",
                     5662 => "00001001",
                     5663 => "00001001",
                     5664 => "11111111",
                     5665 => "11111111",
                     5666 => "00000000",
                     5667 => "00000000",
                     5668 => "00000000",
                     5669 => "00000000",
                     5670 => "00000000",
                     5671 => "00000000",
                     5672 => "11111111",
                     5673 => "00000000",
                     5674 => "11111111",
                     5675 => "11111111",
                     5676 => "11111111",
                     5677 => "11111111",
                     5678 => "11111111",
                     5679 => "11111111",
                     5680 => "11111111",
                     5681 => "11111111",
                     5682 => "00000001",
                     5683 => "01010111",
                     5684 => "00101111",
                     5685 => "01010111",
                     5686 => "00101111",
                     5687 => "01010111",
                     5688 => "11111111",
                     5689 => "00000001",
                     5690 => "11111111",
                     5691 => "10101001",
                     5692 => "11010001",
                     5693 => "10101001",
                     5694 => "11010001",
                     5695 => "10101001",
                     5696 => "11110011",
                     5697 => "11110011",
                     5698 => "11110011",
                     5699 => "11110011",
                     5700 => "11110011",
                     5701 => "11110011",
                     5702 => "11111111",
                     5703 => "00111111",
                     5704 => "10001100",
                     5705 => "10001100",
                     5706 => "10001100",
                     5707 => "10001100",
                     5708 => "10001100",
                     5709 => "10001100",
                     5710 => "11111111",
                     5711 => "00111111",
                     5712 => "11110110",
                     5713 => "11110110",
                     5714 => "11110110",
                     5715 => "11110110",
                     5716 => "11110110",
                     5717 => "11110110",
                     5718 => "11111111",
                     5719 => "11111111",
                     5720 => "00001001",
                     5721 => "00001001",
                     5722 => "00001001",
                     5723 => "00001001",
                     5724 => "00001001",
                     5725 => "00001001",
                     5726 => "11111111",
                     5727 => "11111111",
                     5728 => "00000000",
                     5729 => "00000000",
                     5730 => "00000000",
                     5731 => "00000000",
                     5732 => "00000000",
                     5733 => "00000000",
                     5734 => "11111111",
                     5735 => "11111111",
                     5736 => "11111111",
                     5737 => "11111111",
                     5738 => "11111111",
                     5739 => "11111111",
                     5740 => "11111111",
                     5741 => "11111111",
                     5742 => "11111111",
                     5743 => "11111111",
                     5744 => "00101111",
                     5745 => "01010111",
                     5746 => "00101111",
                     5747 => "01010111",
                     5748 => "00101111",
                     5749 => "01010111",
                     5750 => "11111111",
                     5751 => "11111100",
                     5752 => "11010001",
                     5753 => "10101001",
                     5754 => "11010001",
                     5755 => "10101001",
                     5756 => "11010001",
                     5757 => "10101001",
                     5758 => "11111111",
                     5759 => "11111100",
                     5760 => "00111100",
                     5761 => "00111100",
                     5762 => "00111100",
                     5763 => "00111100",
                     5764 => "00111100",
                     5765 => "00111100",
                     5766 => "00111100",
                     5767 => "00111100",
                     5768 => "00100011",
                     5769 => "00100011",
                     5770 => "00100011",
                     5771 => "00100011",
                     5772 => "00100011",
                     5773 => "00100011",
                     5774 => "00100011",
                     5775 => "00100011",
                     5776 => "11111011",
                     5777 => "11111011",
                     5778 => "11111011",
                     5779 => "11111011",
                     5780 => "11111011",
                     5781 => "11111011",
                     5782 => "11111011",
                     5783 => "11111011",
                     5784 => "00000100",
                     5785 => "00000100",
                     5786 => "00000100",
                     5787 => "00000100",
                     5788 => "00000100",
                     5789 => "00000100",
                     5790 => "00000100",
                     5791 => "00000100",
                     5792 => "10111100",
                     5793 => "01011100",
                     5794 => "10111100",
                     5795 => "01011100",
                     5796 => "10111100",
                     5797 => "01011100",
                     5798 => "10111100",
                     5799 => "01011100",
                     5800 => "01000100",
                     5801 => "10100100",
                     5802 => "01000100",
                     5803 => "10100100",
                     5804 => "01000100",
                     5805 => "10100100",
                     5806 => "01000100",
                     5807 => "10100100",
                     5808 => "00011111",
                     5809 => "00100000",
                     5810 => "01000000",
                     5811 => "01000000",
                     5812 => "10000000",
                     5813 => "10000000",
                     5814 => "10000000",
                     5815 => "10000001",
                     5816 => "00011111",
                     5817 => "00111111",
                     5818 => "01111111",
                     5819 => "01111111",
                     5820 => "11111111",
                     5821 => "11111111",
                     5822 => "11111111",
                     5823 => "11111110",
                     5824 => "11111111",
                     5825 => "10000000",
                     5826 => "10000000",
                     5827 => "11000000",
                     5828 => "11111111",
                     5829 => "11111111",
                     5830 => "11111110",
                     5831 => "11111110",
                     5832 => "11111111",
                     5833 => "01111111",
                     5834 => "01111111",
                     5835 => "00111111",
                     5836 => "00000000",
                     5837 => "00000000",
                     5838 => "00000001",
                     5839 => "00000001",
                     5840 => "11111111",
                     5841 => "01111111",
                     5842 => "01111111",
                     5843 => "11111111",
                     5844 => "11111111",
                     5845 => "00000111",
                     5846 => "00000011",
                     5847 => "00000011",
                     5848 => "11111111",
                     5849 => "10000000",
                     5850 => "10000000",
                     5851 => "00000000",
                     5852 => "00000000",
                     5853 => "11111000",
                     5854 => "11111100",
                     5855 => "11111100",
                     5856 => "11111111",
                     5857 => "00000000",
                     5858 => "00000000",
                     5859 => "00000000",
                     5860 => "00000000",
                     5861 => "10000001",
                     5862 => "11000011",
                     5863 => "11111111",
                     5864 => "11111111",
                     5865 => "11111111",
                     5866 => "11111111",
                     5867 => "11111111",
                     5868 => "11111111",
                     5869 => "01111110",
                     5870 => "00111100",
                     5871 => "00000000",
                     5872 => "11111000",
                     5873 => "11111100",
                     5874 => "11111110",
                     5875 => "11111110",
                     5876 => "11100011",
                     5877 => "11000001",
                     5878 => "10000001",
                     5879 => "10000001",
                     5880 => "11111000",
                     5881 => "00000100",
                     5882 => "00000010",
                     5883 => "00000010",
                     5884 => "00011101",
                     5885 => "00111111",
                     5886 => "01111111",
                     5887 => "01111111",
                     5888 => "10000011",
                     5889 => "11111111",
                     5890 => "11111111",
                     5891 => "11111111",
                     5892 => "11111111",
                     5893 => "11111111",
                     5894 => "01111111",
                     5895 => "00011111",
                     5896 => "11111100",
                     5897 => "10000000",
                     5898 => "10000000",
                     5899 => "10000000",
                     5900 => "10000000",
                     5901 => "10000000",
                     5902 => "01100000",
                     5903 => "00011111",
                     5904 => "11111100",
                     5905 => "11111100",
                     5906 => "11111100",
                     5907 => "11111100",
                     5908 => "11111110",
                     5909 => "11111110",
                     5910 => "11111111",
                     5911 => "11111111",
                     5912 => "00000011",
                     5913 => "00000011",
                     5914 => "00000011",
                     5915 => "00000011",
                     5916 => "00000001",
                     5917 => "00000001",
                     5918 => "00000000",
                     5919 => "11111111",
                     5920 => "00000001",
                     5921 => "00000001",
                     5922 => "00000001",
                     5923 => "00000001",
                     5924 => "00000011",
                     5925 => "00000011",
                     5926 => "00000111",
                     5927 => "11111111",
                     5928 => "11111110",
                     5929 => "11111110",
                     5930 => "11111110",
                     5931 => "11111110",
                     5932 => "11111100",
                     5933 => "11111100",
                     5934 => "11111000",
                     5935 => "11111111",
                     5936 => "11111111",
                     5937 => "11111111",
                     5938 => "11111111",
                     5939 => "11111111",
                     5940 => "11111111",
                     5941 => "11111111",
                     5942 => "11111111",
                     5943 => "11111111",
                     5944 => "00000000",
                     5945 => "00000000",
                     5946 => "00000000",
                     5947 => "00000000",
                     5948 => "00000000",
                     5949 => "00000000",
                     5950 => "00000000",
                     5951 => "11111111",
                     5952 => "10000001",
                     5953 => "11000001",
                     5954 => "11100011",
                     5955 => "11111111",
                     5956 => "11111111",
                     5957 => "11111111",
                     5958 => "11111111",
                     5959 => "11111110",
                     5960 => "01111111",
                     5961 => "00111111",
                     5962 => "00011101",
                     5963 => "00000001",
                     5964 => "00000001",
                     5965 => "00000001",
                     5966 => "00000011",
                     5967 => "11111110",
                     5968 => "11111111",
                     5969 => "11111111",
                     5970 => "11111111",
                     5971 => "11111111",
                     5972 => "11111111",
                     5973 => "11111011",
                     5974 => "10110101",
                     5975 => "11001110",
                     5976 => "10000000",
                     5977 => "10000000",
                     5978 => "10000000",
                     5979 => "10000000",
                     5980 => "10000000",
                     5981 => "10000100",
                     5982 => "11001010",
                     5983 => "10110001",
                     5984 => "11111111",
                     5985 => "11111111",
                     5986 => "11111111",
                     5987 => "11111111",
                     5988 => "11111111",
                     5989 => "11011111",
                     5990 => "10101101",
                     5991 => "01110011",
                     5992 => "00000001",
                     5993 => "00000001",
                     5994 => "00000001",
                     5995 => "00000001",
                     5996 => "00000001",
                     5997 => "00100001",
                     5998 => "01010011",
                     5999 => "10001101",
                     6000 => "01110111",
                     6001 => "01110111",
                     6002 => "01110111",
                     6003 => "01110111",
                     6004 => "01110111",
                     6005 => "01110111",
                     6006 => "01110111",
                     6007 => "01110111",
                     6008 => "00000000",
                     6009 => "00000000",
                     6010 => "00000000",
                     6011 => "00000000",
                     6012 => "01110111",
                     6013 => "11111111",
                     6014 => "11111111",
                     6015 => "11111111",
                     6016 => "00000000",
                     6017 => "00000000",
                     6018 => "00000000",
                     6019 => "00000000",
                     6020 => "00000000",
                     6021 => "00000000",
                     6022 => "00000000",
                     6023 => "11111111",
                     6024 => "11111111",
                     6025 => "11111111",
                     6026 => "11111111",
                     6027 => "11111111",
                     6028 => "11111111",
                     6029 => "11111111",
                     6030 => "11111111",
                     6031 => "11111111",
                     6032 => "01110111",
                     6033 => "01110111",
                     6034 => "01110111",
                     6035 => "01110111",
                     6036 => "00000000",
                     6037 => "00000000",
                     6038 => "00000000",
                     6039 => "00000000",
                     6040 => "11111111",
                     6041 => "11111111",
                     6042 => "11111111",
                     6043 => "01110111",
                     6044 => "01110111",
                     6045 => "01110111",
                     6046 => "01110111",
                     6047 => "01110111",
                     6048 => "00000001",
                     6049 => "00000001",
                     6050 => "00000001",
                     6051 => "00011001",
                     6052 => "00011101",
                     6053 => "00001101",
                     6054 => "00000001",
                     6055 => "11111110",
                     6056 => "11111111",
                     6057 => "11111111",
                     6058 => "11111111",
                     6059 => "11100111",
                     6060 => "11100111",
                     6061 => "11111111",
                     6062 => "11111111",
                     6063 => "11111110",
                     6064 => "00100000",
                     6065 => "01111000",
                     6066 => "01111111",
                     6067 => "11111110",
                     6068 => "11111110",
                     6069 => "11111110",
                     6070 => "11111110",
                     6071 => "11111110",
                     6072 => "00000000",
                     6073 => "00100001",
                     6074 => "00100001",
                     6075 => "01000001",
                     6076 => "01000001",
                     6077 => "01000001",
                     6078 => "01000001",
                     6079 => "01000001",
                     6080 => "00000100",
                     6081 => "10011010",
                     6082 => "11111010",
                     6083 => "11111101",
                     6084 => "11111101",
                     6085 => "11111101",
                     6086 => "11111101",
                     6087 => "11111101",
                     6088 => "00000000",
                     6089 => "10000000",
                     6090 => "10000000",
                     6091 => "10000000",
                     6092 => "10000000",
                     6093 => "10000000",
                     6094 => "10000000",
                     6095 => "10000000",
                     6096 => "01111110",
                     6097 => "00111000",
                     6098 => "00100001",
                     6099 => "00000000",
                     6100 => "00000001",
                     6101 => "00000000",
                     6102 => "00000001",
                     6103 => "00000000",
                     6104 => "00100001",
                     6105 => "00100001",
                     6106 => "00000001",
                     6107 => "00000001",
                     6108 => "00000001",
                     6109 => "00000001",
                     6110 => "00000001",
                     6111 => "00000001",
                     6112 => "11111010",
                     6113 => "10001010",
                     6114 => "10000100",
                     6115 => "10000000",
                     6116 => "10000000",
                     6117 => "10000000",
                     6118 => "10000000",
                     6119 => "10000000",
                     6120 => "10000000",
                     6121 => "10000000",
                     6122 => "10000000",
                     6123 => "10000000",
                     6124 => "10000000",
                     6125 => "10000000",
                     6126 => "10000000",
                     6127 => "10000000",
                     6128 => "00000010",
                     6129 => "00000100",
                     6130 => "00000000",
                     6131 => "00010000",
                     6132 => "00000000",
                     6133 => "01000000",
                     6134 => "10000000",
                     6135 => "00000000",
                     6136 => "00000001",
                     6137 => "00000001",
                     6138 => "00000110",
                     6139 => "00001000",
                     6140 => "00011000",
                     6141 => "00100000",
                     6142 => "00100000",
                     6143 => "11000000",
                     6144 => "00001011",
                     6145 => "00001011",
                     6146 => "00111011",
                     6147 => "00001011",
                     6148 => "11111011",
                     6149 => "00001011",
                     6150 => "00001011",
                     6151 => "00001010",
                     6152 => "00000100",
                     6153 => "00000100",
                     6154 => "11000100",
                     6155 => "11110100",
                     6156 => "11110100",
                     6157 => "00000100",
                     6158 => "00000100",
                     6159 => "00000101",
                     6160 => "10010000",
                     6161 => "00010000",
                     6162 => "00011111",
                     6163 => "00010000",
                     6164 => "00011111",
                     6165 => "00010000",
                     6166 => "00010000",
                     6167 => "10010000",
                     6168 => "01110000",
                     6169 => "11110000",
                     6170 => "11110000",
                     6171 => "11111111",
                     6172 => "11111111",
                     6173 => "11110000",
                     6174 => "11110000",
                     6175 => "01110000",
                     6176 => "00111111",
                     6177 => "01111000",
                     6178 => "11100111",
                     6179 => "11001111",
                     6180 => "01011000",
                     6181 => "01011000",
                     6182 => "01010000",
                     6183 => "10010000",
                     6184 => "11000000",
                     6185 => "10000111",
                     6186 => "00011000",
                     6187 => "10110000",
                     6188 => "11100111",
                     6189 => "11100111",
                     6190 => "11101111",
                     6191 => "11101111",
                     6192 => "10110000",
                     6193 => "11111100",
                     6194 => "11100010",
                     6195 => "11000001",
                     6196 => "11000001",
                     6197 => "10000011",
                     6198 => "10001111",
                     6199 => "01111110",
                     6200 => "01101111",
                     6201 => "01000011",
                     6202 => "01011101",
                     6203 => "00111111",
                     6204 => "00111111",
                     6205 => "01111111",
                     6206 => "01111111",
                     6207 => "11111111",
                     6208 => "11111110",
                     6209 => "00000011",
                     6210 => "00001111",
                     6211 => "10010001",
                     6212 => "01110000",
                     6213 => "01100000",
                     6214 => "00100000",
                     6215 => "00110001",
                     6216 => "00000011",
                     6217 => "11111111",
                     6218 => "11110001",
                     6219 => "01101110",
                     6220 => "11001111",
                     6221 => "11011111",
                     6222 => "11111111",
                     6223 => "11111111",
                     6224 => "00111111",
                     6225 => "00111111",
                     6226 => "00011101",
                     6227 => "00111001",
                     6228 => "01111011",
                     6229 => "11110011",
                     6230 => "10000110",
                     6231 => "11111110",
                     6232 => "11111101",
                     6233 => "11111011",
                     6234 => "11111011",
                     6235 => "11110111",
                     6236 => "11110111",
                     6237 => "00001111",
                     6238 => "01111111",
                     6239 => "11111111",
                     6240 => "11111111",
                     6241 => "11111111",
                     6242 => "11111111",
                     6243 => "11111111",
                     6244 => "11111111",
                     6245 => "10000000",
                     6246 => "10000000",
                     6247 => "11111111",
                     6248 => "11111111",
                     6249 => "10000000",
                     6250 => "10000000",
                     6251 => "10000000",
                     6252 => "10000000",
                     6253 => "11111111",
                     6254 => "11111111",
                     6255 => "10000000",
                     6256 => "11111110",
                     6257 => "11111111",
                     6258 => "11111111",
                     6259 => "11111111",
                     6260 => "11111111",
                     6261 => "00000011",
                     6262 => "00000011",
                     6263 => "11111111",
                     6264 => "11111110",
                     6265 => "00000011",
                     6266 => "00000011",
                     6267 => "00000011",
                     6268 => "00000011",
                     6269 => "11111111",
                     6270 => "11111111",
                     6271 => "00000011",
                     6272 => "00000000",
                     6273 => "11111111",
                     6274 => "11111111",
                     6275 => "11111111",
                     6276 => "11111111",
                     6277 => "11111111",
                     6278 => "00000000",
                     6279 => "00000000",
                     6280 => "00000000",
                     6281 => "11111111",
                     6282 => "00000000",
                     6283 => "00000000",
                     6284 => "00000000",
                     6285 => "00000000",
                     6286 => "11111111",
                     6287 => "11111111",
                     6288 => "00111100",
                     6289 => "11111100",
                     6290 => "11111100",
                     6291 => "11111100",
                     6292 => "11111100",
                     6293 => "11111100",
                     6294 => "00000100",
                     6295 => "00000100",
                     6296 => "00100011",
                     6297 => "11110011",
                     6298 => "00001011",
                     6299 => "00001011",
                     6300 => "00001011",
                     6301 => "00000111",
                     6302 => "11111111",
                     6303 => "11111111",
                     6304 => "11111111",
                     6305 => "11111111",
                     6306 => "11111111",
                     6307 => "11111111",
                     6308 => "10000000",
                     6309 => "11111111",
                     6310 => "11111111",
                     6311 => "11111111",
                     6312 => "10000000",
                     6313 => "10000000",
                     6314 => "10000000",
                     6315 => "10000000",
                     6316 => "11111111",
                     6317 => "10000000",
                     6318 => "10000000",
                     6319 => "10000000",
                     6320 => "11111111",
                     6321 => "11111111",
                     6322 => "11111111",
                     6323 => "11111111",
                     6324 => "00000011",
                     6325 => "11111111",
                     6326 => "11111111",
                     6327 => "11111111",
                     6328 => "00000011",
                     6329 => "00000011",
                     6330 => "00000011",
                     6331 => "00000011",
                     6332 => "11111111",
                     6333 => "00000011",
                     6334 => "00000011",
                     6335 => "00000011",
                     6336 => "11111111",
                     6337 => "11111111",
                     6338 => "11111111",
                     6339 => "11111111",
                     6340 => "11111111",
                     6341 => "00000000",
                     6342 => "11111111",
                     6343 => "11111111",
                     6344 => "00000000",
                     6345 => "00000000",
                     6346 => "00000000",
                     6347 => "00000000",
                     6348 => "00000000",
                     6349 => "11111111",
                     6350 => "00000000",
                     6351 => "00000000",
                     6352 => "11111100",
                     6353 => "11111100",
                     6354 => "11111110",
                     6355 => "11111110",
                     6356 => "11111110",
                     6357 => "00000010",
                     6358 => "11111110",
                     6359 => "11111110",
                     6360 => "00000111",
                     6361 => "00000111",
                     6362 => "00000011",
                     6363 => "00000011",
                     6364 => "00000011",
                     6365 => "11111111",
                     6366 => "00000011",
                     6367 => "00000011",
                     6368 => "11111111",
                     6369 => "10000000",
                     6370 => "10000000",
                     6371 => "10000000",
                     6372 => "10000000",
                     6373 => "10000000",
                     6374 => "10000000",
                     6375 => "10000000",
                     6376 => "10000000",
                     6377 => "11111111",
                     6378 => "11111111",
                     6379 => "11111111",
                     6380 => "11111111",
                     6381 => "11111111",
                     6382 => "11111111",
                     6383 => "11111111",
                     6384 => "11111111",
                     6385 => "00000011",
                     6386 => "00000011",
                     6387 => "00000011",
                     6388 => "00000011",
                     6389 => "00000011",
                     6390 => "00000011",
                     6391 => "00000011",
                     6392 => "00000011",
                     6393 => "11111111",
                     6394 => "11111111",
                     6395 => "11111111",
                     6396 => "11111111",
                     6397 => "11111111",
                     6398 => "11111111",
                     6399 => "11111111",
                     6400 => "00000010",
                     6401 => "00000010",
                     6402 => "00000010",
                     6403 => "00000010",
                     6404 => "00000010",
                     6405 => "00000010",
                     6406 => "00000100",
                     6407 => "00000100",
                     6408 => "11111111",
                     6409 => "11111111",
                     6410 => "11111111",
                     6411 => "11111111",
                     6412 => "11111111",
                     6413 => "11111111",
                     6414 => "11111111",
                     6415 => "11111111",
                     6416 => "10000000",
                     6417 => "10000000",
                     6418 => "10101010",
                     6419 => "11010101",
                     6420 => "10101010",
                     6421 => "11111111",
                     6422 => "11111111",
                     6423 => "11111111",
                     6424 => "11111111",
                     6425 => "11111111",
                     6426 => "11010101",
                     6427 => "10101010",
                     6428 => "11010101",
                     6429 => "10000000",
                     6430 => "10000000",
                     6431 => "11111111",
                     6432 => "00000011",
                     6433 => "00000011",
                     6434 => "10101011",
                     6435 => "01010111",
                     6436 => "10101011",
                     6437 => "11111111",
                     6438 => "11111111",
                     6439 => "11111110",
                     6440 => "11111111",
                     6441 => "11111111",
                     6442 => "01010111",
                     6443 => "10101011",
                     6444 => "01010111",
                     6445 => "00000011",
                     6446 => "00000011",
                     6447 => "11111110",
                     6448 => "00000000",
                     6449 => "01010101",
                     6450 => "10101010",
                     6451 => "01010101",
                     6452 => "11111111",
                     6453 => "11111111",
                     6454 => "11111111",
                     6455 => "00000000",
                     6456 => "11111111",
                     6457 => "10101010",
                     6458 => "01010101",
                     6459 => "10101010",
                     6460 => "00000000",
                     6461 => "00000000",
                     6462 => "11111111",
                     6463 => "00000000",
                     6464 => "00000100",
                     6465 => "01010100",
                     6466 => "10101100",
                     6467 => "01011100",
                     6468 => "11111100",
                     6469 => "11111100",
                     6470 => "11111100",
                     6471 => "00111100",
                     6472 => "11111111",
                     6473 => "10101111",
                     6474 => "01010111",
                     6475 => "10101011",
                     6476 => "00001011",
                     6477 => "00001011",
                     6478 => "11110011",
                     6479 => "00100011",
                     6480 => "00111111",
                     6481 => "00111111",
                     6482 => "00111111",
                     6483 => "00111111",
                     6484 => "00000000",
                     6485 => "00000000",
                     6486 => "00000000",
                     6487 => "11111111",
                     6488 => "11111111",
                     6489 => "11111111",
                     6490 => "11111111",
                     6491 => "11111111",
                     6492 => "11111111",
                     6493 => "11111111",
                     6494 => "11111111",
                     6495 => "11111111",
                     6496 => "01111110",
                     6497 => "01111100",
                     6498 => "01111100",
                     6499 => "01111000",
                     6500 => "00000000",
                     6501 => "00000000",
                     6502 => "00000000",
                     6503 => "11111111",
                     6504 => "11111111",
                     6505 => "11111111",
                     6506 => "11111111",
                     6507 => "11111111",
                     6508 => "11111111",
                     6509 => "11111111",
                     6510 => "11111111",
                     6511 => "11111111",
                     6512 => "00011111",
                     6513 => "00001111",
                     6514 => "00001111",
                     6515 => "00000111",
                     6516 => "00000000",
                     6517 => "00000000",
                     6518 => "00000000",
                     6519 => "11111111",
                     6520 => "11111111",
                     6521 => "11111111",
                     6522 => "11111111",
                     6523 => "11111111",
                     6524 => "11111111",
                     6525 => "11111111",
                     6526 => "11111111",
                     6527 => "11111111",
                     6528 => "11111110",
                     6529 => "11111100",
                     6530 => "11111100",
                     6531 => "11111000",
                     6532 => "00000000",
                     6533 => "00000000",
                     6534 => "00000000",
                     6535 => "11111111",
                     6536 => "11111111",
                     6537 => "11111111",
                     6538 => "11111111",
                     6539 => "11111111",
                     6540 => "11111111",
                     6541 => "11111111",
                     6542 => "11111111",
                     6543 => "11111111",
                     6544 => "00000000",
                     6545 => "00000000",
                     6546 => "00000000",
                     6547 => "00000000",
                     6548 => "11111111",
                     6549 => "11111111",
                     6550 => "00000000",
                     6551 => "00000000",
                     6552 => "00000000",
                     6553 => "00000000",
                     6554 => "00000000",
                     6555 => "00000000",
                     6556 => "00000000",
                     6557 => "00000000",
                     6558 => "00000000",
                     6559 => "00000000",
                     6560 => "00011000",
                     6561 => "00011000",
                     6562 => "00011000",
                     6563 => "00011000",
                     6564 => "00011000",
                     6565 => "00011000",
                     6566 => "00011000",
                     6567 => "00011000",
                     6568 => "00000000",
                     6569 => "00000000",
                     6570 => "00000000",
                     6571 => "00000000",
                     6572 => "00000000",
                     6573 => "00000000",
                     6574 => "00000000",
                     6575 => "00000000",
                     6576 => "00000111",
                     6577 => "00011111",
                     6578 => "00111111",
                     6579 => "11111111",
                     6580 => "01111111",
                     6581 => "01111111",
                     6582 => "11111111",
                     6583 => "11111111",
                     6584 => "11111111",
                     6585 => "11111111",
                     6586 => "11111111",
                     6587 => "11111111",
                     6588 => "11111111",
                     6589 => "11111111",
                     6590 => "11111111",
                     6591 => "11111111",
                     6592 => "11100001",
                     6593 => "11111001",
                     6594 => "11111101",
                     6595 => "11111111",
                     6596 => "11111110",
                     6597 => "11111110",
                     6598 => "11111111",
                     6599 => "11111111",
                     6600 => "11111111",
                     6601 => "11111111",
                     6602 => "11111111",
                     6603 => "11111111",
                     6604 => "11111111",
                     6605 => "11111111",
                     6606 => "11111111",
                     6607 => "11111111",
                     6608 => "11110000",
                     6609 => "00010000",
                     6610 => "00010000",
                     6611 => "00010000",
                     6612 => "00010000",
                     6613 => "00010000",
                     6614 => "00010000",
                     6615 => "11111111",
                     6616 => "00000000",
                     6617 => "11100000",
                     6618 => "11100000",
                     6619 => "11100000",
                     6620 => "11100000",
                     6621 => "11100000",
                     6622 => "11100000",
                     6623 => "11100000",
                     6624 => "00011111",
                     6625 => "00010000",
                     6626 => "00010000",
                     6627 => "00010000",
                     6628 => "00010000",
                     6629 => "00010000",
                     6630 => "00010000",
                     6631 => "11111111",
                     6632 => "00000000",
                     6633 => "00001111",
                     6634 => "00001111",
                     6635 => "00001111",
                     6636 => "00001111",
                     6637 => "00001111",
                     6638 => "00001111",
                     6639 => "00001111",
                     6640 => "10010010",
                     6641 => "10010010",
                     6642 => "10010010",
                     6643 => "11111110",
                     6644 => "11111110",
                     6645 => "00000000",
                     6646 => "00000000",
                     6647 => "00000000",
                     6648 => "01001000",
                     6649 => "01001000",
                     6650 => "01101100",
                     6651 => "00000000",
                     6652 => "00000000",
                     6653 => "00000000",
                     6654 => "11111110",
                     6655 => "00000000",
                     6656 => "00001010",
                     6657 => "00001010",
                     6658 => "00111010",
                     6659 => "00001010",
                     6660 => "11111011",
                     6661 => "00001011",
                     6662 => "00001011",
                     6663 => "00001011",
                     6664 => "00000101",
                     6665 => "00000101",
                     6666 => "11000101",
                     6667 => "11110101",
                     6668 => "11110100",
                     6669 => "00000100",
                     6670 => "00000100",
                     6671 => "00000100",
                     6672 => "10010000",
                     6673 => "10010000",
                     6674 => "10011111",
                     6675 => "10010000",
                     6676 => "10011111",
                     6677 => "10010000",
                     6678 => "10010000",
                     6679 => "10010000",
                     6680 => "01110000",
                     6681 => "01110000",
                     6682 => "01110000",
                     6683 => "01111111",
                     6684 => "01111111",
                     6685 => "01110000",
                     6686 => "01110000",
                     6687 => "01110000",
                     6688 => "00000001",
                     6689 => "00000001",
                     6690 => "00000001",
                     6691 => "00000001",
                     6692 => "00000001",
                     6693 => "00000001",
                     6694 => "00000001",
                     6695 => "00000001",
                     6696 => "00000000",
                     6697 => "00000000",
                     6698 => "00000000",
                     6699 => "00000000",
                     6700 => "00000000",
                     6701 => "00000000",
                     6702 => "00000000",
                     6703 => "00000000",
                     6704 => "10000000",
                     6705 => "10000000",
                     6706 => "10000000",
                     6707 => "10000000",
                     6708 => "10000000",
                     6709 => "10000000",
                     6710 => "10000000",
                     6711 => "10000000",
                     6712 => "00000000",
                     6713 => "00000000",
                     6714 => "00000000",
                     6715 => "00000000",
                     6716 => "00000000",
                     6717 => "00000000",
                     6718 => "00000000",
                     6719 => "00000000",
                     6720 => "00001000",
                     6721 => "10001000",
                     6722 => "10010001",
                     6723 => "11010001",
                     6724 => "01010011",
                     6725 => "01010011",
                     6726 => "01110011",
                     6727 => "00111111",
                     6728 => "11111111",
                     6729 => "11111111",
                     6730 => "11111111",
                     6731 => "11111111",
                     6732 => "11111111",
                     6733 => "11111110",
                     6734 => "10111110",
                     6735 => "11001110",
                     6736 => "00000000",
                     6737 => "00000000",
                     6738 => "00000111",
                     6739 => "00001111",
                     6740 => "00001100",
                     6741 => "00011011",
                     6742 => "00011011",
                     6743 => "00011011",
                     6744 => "00000000",
                     6745 => "00000000",
                     6746 => "00000000",
                     6747 => "00000000",
                     6748 => "00000011",
                     6749 => "00000100",
                     6750 => "00000100",
                     6751 => "00000100",
                     6752 => "00000000",
                     6753 => "00000000",
                     6754 => "11100000",
                     6755 => "11110000",
                     6756 => "11110000",
                     6757 => "11111000",
                     6758 => "11111000",
                     6759 => "11111000",
                     6760 => "00000000",
                     6761 => "00000000",
                     6762 => "01100000",
                     6763 => "00110000",
                     6764 => "00110000",
                     6765 => "10011000",
                     6766 => "10011000",
                     6767 => "10011000",
                     6768 => "00011011",
                     6769 => "00011011",
                     6770 => "00011011",
                     6771 => "00011011",
                     6772 => "00011011",
                     6773 => "00001111",
                     6774 => "00001111",
                     6775 => "00000111",
                     6776 => "00000100",
                     6777 => "00000100",
                     6778 => "00000100",
                     6779 => "00000100",
                     6780 => "00000100",
                     6781 => "00000011",
                     6782 => "00000000",
                     6783 => "00000000",
                     6784 => "11111000",
                     6785 => "11111000",
                     6786 => "11111000",
                     6787 => "11111000",
                     6788 => "11111000",
                     6789 => "11110000",
                     6790 => "11110000",
                     6791 => "11100000",
                     6792 => "10011000",
                     6793 => "10011000",
                     6794 => "10011000",
                     6795 => "10011000",
                     6796 => "10011000",
                     6797 => "00110000",
                     6798 => "00110000",
                     6799 => "01100000",
                     6800 => "11110001",
                     6801 => "00010001",
                     6802 => "00010001",
                     6803 => "00011111",
                     6804 => "00010000",
                     6805 => "00010000",
                     6806 => "00010000",
                     6807 => "11111111",
                     6808 => "00001111",
                     6809 => "11101111",
                     6810 => "11101111",
                     6811 => "11101111",
                     6812 => "11101111",
                     6813 => "11101111",
                     6814 => "11101111",
                     6815 => "11100000",
                     6816 => "00011111",
                     6817 => "00010000",
                     6818 => "00010000",
                     6819 => "11110000",
                     6820 => "00010000",
                     6821 => "00010000",
                     6822 => "00010000",
                     6823 => "11111111",
                     6824 => "11100000",
                     6825 => "11101111",
                     6826 => "11101111",
                     6827 => "11101111",
                     6828 => "11101111",
                     6829 => "11101111",
                     6830 => "11101111",
                     6831 => "00001111",
                     6832 => "01111111",
                     6833 => "10111111",
                     6834 => "11011111",
                     6835 => "11101111",
                     6836 => "11110000",
                     6837 => "11110000",
                     6838 => "11110000",
                     6839 => "11110000",
                     6840 => "10000000",
                     6841 => "01000000",
                     6842 => "00100000",
                     6843 => "00010000",
                     6844 => "00001111",
                     6845 => "00001111",
                     6846 => "00001111",
                     6847 => "00001111",
                     6848 => "11110000",
                     6849 => "11110000",
                     6850 => "11110000",
                     6851 => "11110000",
                     6852 => "11111111",
                     6853 => "11111111",
                     6854 => "11111111",
                     6855 => "11111111",
                     6856 => "00001111",
                     6857 => "00001111",
                     6858 => "00001111",
                     6859 => "00001111",
                     6860 => "00011111",
                     6861 => "00111111",
                     6862 => "01111111",
                     6863 => "11111111",
                     6864 => "11111111",
                     6865 => "11111111",
                     6866 => "11111111",
                     6867 => "11111111",
                     6868 => "00001111",
                     6869 => "00001111",
                     6870 => "00001111",
                     6871 => "00001111",
                     6872 => "00000001",
                     6873 => "00000011",
                     6874 => "00000111",
                     6875 => "00001111",
                     6876 => "11111111",
                     6877 => "11111111",
                     6878 => "11111111",
                     6879 => "11111111",
                     6880 => "00001111",
                     6881 => "00001111",
                     6882 => "00001111",
                     6883 => "00001111",
                     6884 => "11110111",
                     6885 => "11111011",
                     6886 => "11111101",
                     6887 => "11111110",
                     6888 => "11111111",
                     6889 => "11111111",
                     6890 => "11111111",
                     6891 => "11111111",
                     6892 => "11111111",
                     6893 => "11111111",
                     6894 => "11111111",
                     6895 => "11111111",
                     6896 => "00000000",
                     6897 => "00000000",
                     6898 => "00000000",
                     6899 => "00000000",
                     6900 => "00000000",
                     6901 => "00000000",
                     6902 => "00011000",
                     6903 => "00011000",
                     6904 => "00000000",
                     6905 => "00000000",
                     6906 => "00000000",
                     6907 => "00000000",
                     6908 => "00000000",
                     6909 => "00000000",
                     6910 => "00000000",
                     6911 => "00000000",
                     6912 => "00011111",
                     6913 => "00111111",
                     6914 => "01111111",
                     6915 => "01111111",
                     6916 => "01111111",
                     6917 => "11111111",
                     6918 => "11111111",
                     6919 => "11111111",
                     6920 => "00011111",
                     6921 => "00100000",
                     6922 => "01000000",
                     6923 => "01000000",
                     6924 => "01000000",
                     6925 => "10000000",
                     6926 => "10000010",
                     6927 => "10000010",
                     6928 => "11111111",
                     6929 => "11111111",
                     6930 => "11111111",
                     6931 => "01111111",
                     6932 => "01111111",
                     6933 => "01111111",
                     6934 => "00111111",
                     6935 => "00011110",
                     6936 => "10000010",
                     6937 => "10000000",
                     6938 => "10100000",
                     6939 => "01000100",
                     6940 => "01000011",
                     6941 => "01000000",
                     6942 => "00100001",
                     6943 => "00011110",
                     6944 => "11111000",
                     6945 => "11111100",
                     6946 => "11111110",
                     6947 => "11111110",
                     6948 => "11111110",
                     6949 => "11111111",
                     6950 => "11111111",
                     6951 => "11111111",
                     6952 => "11111000",
                     6953 => "00000100",
                     6954 => "00000010",
                     6955 => "00000010",
                     6956 => "00000010",
                     6957 => "00000001",
                     6958 => "01000001",
                     6959 => "01000001",
                     6960 => "11111111",
                     6961 => "11111111",
                     6962 => "11111111",
                     6963 => "11111110",
                     6964 => "11111110",
                     6965 => "11111110",
                     6966 => "11111100",
                     6967 => "01111000",
                     6968 => "01000001",
                     6969 => "00000001",
                     6970 => "00000101",
                     6971 => "00100010",
                     6972 => "11000010",
                     6973 => "00000010",
                     6974 => "10000100",
                     6975 => "01111000",
                     6976 => "01111111",
                     6977 => "10000000",
                     6978 => "10000000",
                     6979 => "10000000",
                     6980 => "10000000",
                     6981 => "10000000",
                     6982 => "10000000",
                     6983 => "10000000",
                     6984 => "10000000",
                     6985 => "01111111",
                     6986 => "01111111",
                     6987 => "01111111",
                     6988 => "01111111",
                     6989 => "01111111",
                     6990 => "01111111",
                     6991 => "01111111",
                     6992 => "11011110",
                     6993 => "01100001",
                     6994 => "01100001",
                     6995 => "01100001",
                     6996 => "01110001",
                     6997 => "01011110",
                     6998 => "01111111",
                     6999 => "01100001",
                     7000 => "01100001",
                     7001 => "11011111",
                     7002 => "11011111",
                     7003 => "11011111",
                     7004 => "11011111",
                     7005 => "11111111",
                     7006 => "11000001",
                     7007 => "11011111",
                     7008 => "10000000",
                     7009 => "10000000",
                     7010 => "11000000",
                     7011 => "11110000",
                     7012 => "10111111",
                     7013 => "10001111",
                     7014 => "10000001",
                     7015 => "01111110",
                     7016 => "01111111",
                     7017 => "01111111",
                     7018 => "11111111",
                     7019 => "00111111",
                     7020 => "01001111",
                     7021 => "01110001",
                     7022 => "01111111",
                     7023 => "11111111",
                     7024 => "01100001",
                     7025 => "01100001",
                     7026 => "11000001",
                     7027 => "11000001",
                     7028 => "10000001",
                     7029 => "10000001",
                     7030 => "10000011",
                     7031 => "11111110",
                     7032 => "11011111",
                     7033 => "11011111",
                     7034 => "10111111",
                     7035 => "10111111",
                     7036 => "01111111",
                     7037 => "01111111",
                     7038 => "01111111",
                     7039 => "01111111",
                     7040 => "00000000",
                     7041 => "00000000",
                     7042 => "00000011",
                     7043 => "00001111",
                     7044 => "00011111",
                     7045 => "00111111",
                     7046 => "01111111",
                     7047 => "01111111",
                     7048 => "00000000",
                     7049 => "00000000",
                     7050 => "00000011",
                     7051 => "00001100",
                     7052 => "00010000",
                     7053 => "00100000",
                     7054 => "01000000",
                     7055 => "01000000",
                     7056 => "00000000",
                     7057 => "00000000",
                     7058 => "11000000",
                     7059 => "11110000",
                     7060 => "11111000",
                     7061 => "11111100",
                     7062 => "11111110",
                     7063 => "11111110",
                     7064 => "00000000",
                     7065 => "00000000",
                     7066 => "11000000",
                     7067 => "00110000",
                     7068 => "00001000",
                     7069 => "00000100",
                     7070 => "00000010",
                     7071 => "00000010",
                     7072 => "11111111",
                     7073 => "11111111",
                     7074 => "11111111",
                     7075 => "11111111",
                     7076 => "11111111",
                     7077 => "11111111",
                     7078 => "11111111",
                     7079 => "11111111",
                     7080 => "10000000",
                     7081 => "10000000",
                     7082 => "10000000",
                     7083 => "10000000",
                     7084 => "10000000",
                     7085 => "10000000",
                     7086 => "10000000",
                     7087 => "10000000",
                     7088 => "11111111",
                     7089 => "11111111",
                     7090 => "11111111",
                     7091 => "11111111",
                     7092 => "11111111",
                     7093 => "11111111",
                     7094 => "11111111",
                     7095 => "11111111",
                     7096 => "00000001",
                     7097 => "00000001",
                     7098 => "00000001",
                     7099 => "00000001",
                     7100 => "00000001",
                     7101 => "00000001",
                     7102 => "00000001",
                     7103 => "00000001",
                     7104 => "01111111",
                     7105 => "01111111",
                     7106 => "01111111",
                     7107 => "00111111",
                     7108 => "00111111",
                     7109 => "00011111",
                     7110 => "00001111",
                     7111 => "00000111",
                     7112 => "01000000",
                     7113 => "01000000",
                     7114 => "01000000",
                     7115 => "00100000",
                     7116 => "00110000",
                     7117 => "00011100",
                     7118 => "00001111",
                     7119 => "00000111",
                     7120 => "11111110",
                     7121 => "11111110",
                     7122 => "11111110",
                     7123 => "11111100",
                     7124 => "11111100",
                     7125 => "11111000",
                     7126 => "11110000",
                     7127 => "11110000",
                     7128 => "00000010",
                     7129 => "00000010",
                     7130 => "00000010",
                     7131 => "00000100",
                     7132 => "00001100",
                     7133 => "00111000",
                     7134 => "11110000",
                     7135 => "11110000",
                     7136 => "00001111",
                     7137 => "00001111",
                     7138 => "00001111",
                     7139 => "00001111",
                     7140 => "00001111",
                     7141 => "00001111",
                     7142 => "00000111",
                     7143 => "00001111",
                     7144 => "00001000",
                     7145 => "00001000",
                     7146 => "00001000",
                     7147 => "00001000",
                     7148 => "00001000",
                     7149 => "00001100",
                     7150 => "00000101",
                     7151 => "00001010",
                     7152 => "11110000",
                     7153 => "11110000",
                     7154 => "11110000",
                     7155 => "11110000",
                     7156 => "11110000",
                     7157 => "11110000",
                     7158 => "11100000",
                     7159 => "11110000",
                     7160 => "00010000",
                     7161 => "01010000",
                     7162 => "01010000",
                     7163 => "01010000",
                     7164 => "01010000",
                     7165 => "00110000",
                     7166 => "10100000",
                     7167 => "01010000",
                     7168 => "10000001",
                     7169 => "11000001",
                     7170 => "10100011",
                     7171 => "10100011",
                     7172 => "10011101",
                     7173 => "10000001",
                     7174 => "10000001",
                     7175 => "10000001",
                     7176 => "00000000",
                     7177 => "01000001",
                     7178 => "00100010",
                     7179 => "00100010",
                     7180 => "00011100",
                     7181 => "00000000",
                     7182 => "00000000",
                     7183 => "00000000",
                     7184 => "11100011",
                     7185 => "11110111",
                     7186 => "11000001",
                     7187 => "11000001",
                     7188 => "11000001",
                     7189 => "11000001",
                     7190 => "11110111",
                     7191 => "11100011",
                     7192 => "11100011",
                     7193 => "00010100",
                     7194 => "00111110",
                     7195 => "00111110",
                     7196 => "00111110",
                     7197 => "00111110",
                     7198 => "00010100",
                     7199 => "11100011",
                     7200 => "00000000",
                     7201 => "00000000",
                     7202 => "00000111",
                     7203 => "00001111",
                     7204 => "00001100",
                     7205 => "00011011",
                     7206 => "00011011",
                     7207 => "00011011",
                     7208 => "11111111",
                     7209 => "11111111",
                     7210 => "11111000",
                     7211 => "11110000",
                     7212 => "11110000",
                     7213 => "11100000",
                     7214 => "11100000",
                     7215 => "11100000",
                     7216 => "00000000",
                     7217 => "00000000",
                     7218 => "11100000",
                     7219 => "11110000",
                     7220 => "11110000",
                     7221 => "11111000",
                     7222 => "11111000",
                     7223 => "11111000",
                     7224 => "11111111",
                     7225 => "11111111",
                     7226 => "01111111",
                     7227 => "00111111",
                     7228 => "00111111",
                     7229 => "10011111",
                     7230 => "10011111",
                     7231 => "10011111",
                     7232 => "00011011",
                     7233 => "00011011",
                     7234 => "00011011",
                     7235 => "00011011",
                     7236 => "00011011",
                     7237 => "00001111",
                     7238 => "00001111",
                     7239 => "00000111",
                     7240 => "11100000",
                     7241 => "11100000",
                     7242 => "11100000",
                     7243 => "11100000",
                     7244 => "11100000",
                     7245 => "11110011",
                     7246 => "11110000",
                     7247 => "11111000",
                     7248 => "11111000",
                     7249 => "11111000",
                     7250 => "11111000",
                     7251 => "11111000",
                     7252 => "11111000",
                     7253 => "11110000",
                     7254 => "11110000",
                     7255 => "11100000",
                     7256 => "10011111",
                     7257 => "10011111",
                     7258 => "10011111",
                     7259 => "10011111",
                     7260 => "10011111",
                     7261 => "00111111",
                     7262 => "00111111",
                     7263 => "01111111",
                     7264 => "11100000",
                     7265 => "11111111",
                     7266 => "11111111",
                     7267 => "11111111",
                     7268 => "11111111",
                     7269 => "11111111",
                     7270 => "11111111",
                     7271 => "11111111",
                     7272 => "00000000",
                     7273 => "01110000",
                     7274 => "00011111",
                     7275 => "00010000",
                     7276 => "01110000",
                     7277 => "01111111",
                     7278 => "01111111",
                     7279 => "01111111",
                     7280 => "00000111",
                     7281 => "11111111",
                     7282 => "11111111",
                     7283 => "11111111",
                     7284 => "11111111",
                     7285 => "11111111",
                     7286 => "11111111",
                     7287 => "11111111",
                     7288 => "00000000",
                     7289 => "00000011",
                     7290 => "11111000",
                     7291 => "00000000",
                     7292 => "00000011",
                     7293 => "11111011",
                     7294 => "11111011",
                     7295 => "11111011",
                     7296 => "11111111",
                     7297 => "11111111",
                     7298 => "11111111",
                     7299 => "11111111",
                     7300 => "11111111",
                     7301 => "11111110",
                     7302 => "11111111",
                     7303 => "11101111",
                     7304 => "01111100",
                     7305 => "01111011",
                     7306 => "01110110",
                     7307 => "01110101",
                     7308 => "01110101",
                     7309 => "01110111",
                     7310 => "00010111",
                     7311 => "01100111",
                     7312 => "11111111",
                     7313 => "11011111",
                     7314 => "11101111",
                     7315 => "10101111",
                     7316 => "10101111",
                     7317 => "01101111",
                     7318 => "11101111",
                     7319 => "11100111",
                     7320 => "00111011",
                     7321 => "11111011",
                     7322 => "01111011",
                     7323 => "11111011",
                     7324 => "11111011",
                     7325 => "11110011",
                     7326 => "11111000",
                     7327 => "11110011",
                     7328 => "00011111",
                     7329 => "00011111",
                     7330 => "00111111",
                     7331 => "00111111",
                     7332 => "01110000",
                     7333 => "01100011",
                     7334 => "11100111",
                     7335 => "11100101",
                     7336 => "00001111",
                     7337 => "00001111",
                     7338 => "00011111",
                     7339 => "00011111",
                     7340 => "00111111",
                     7341 => "00111100",
                     7342 => "01111000",
                     7343 => "01111010",
                     7344 => "11110000",
                     7345 => "11110000",
                     7346 => "11111000",
                     7347 => "11111000",
                     7348 => "00001100",
                     7349 => "11000100",
                     7350 => "11100100",
                     7351 => "10100110",
                     7352 => "11111000",
                     7353 => "11111000",
                     7354 => "11111100",
                     7355 => "11111100",
                     7356 => "11111110",
                     7357 => "00111110",
                     7358 => "00011110",
                     7359 => "01011111",
                     7360 => "11101001",
                     7361 => "11101001",
                     7362 => "11101001",
                     7363 => "11101111",
                     7364 => "11100010",
                     7365 => "11100011",
                     7366 => "11110000",
                     7367 => "11111111",
                     7368 => "01110110",
                     7369 => "01110110",
                     7370 => "01110110",
                     7371 => "01110000",
                     7372 => "01111101",
                     7373 => "01111100",
                     7374 => "01111111",
                     7375 => "01111111",
                     7376 => "10010110",
                     7377 => "10010110",
                     7378 => "10010110",
                     7379 => "11110110",
                     7380 => "01000110",
                     7381 => "11000110",
                     7382 => "00001110",
                     7383 => "11111110",
                     7384 => "01101111",
                     7385 => "01101111",
                     7386 => "01101111",
                     7387 => "00001111",
                     7388 => "10111111",
                     7389 => "00111111",
                     7390 => "11111111",
                     7391 => "11111111",
                     7392 => "00000000",
                     7393 => "00000000",
                     7394 => "00000000",
                     7395 => "00000000",
                     7396 => "00000000",
                     7397 => "00000000",
                     7398 => "01111110",
                     7399 => "00111100",
                     7400 => "00111100",
                     7401 => "01111110",
                     7402 => "01111110",
                     7403 => "11111111",
                     7404 => "11111111",
                     7405 => "11111111",
                     7406 => "01000010",
                     7407 => "00000000",
                     7408 => "00111100",
                     7409 => "01000010",
                     7410 => "10011001",
                     7411 => "10100001",
                     7412 => "10100001",
                     7413 => "10011001",
                     7414 => "01000010",
                     7415 => "00111100",
                     7416 => "00000000",
                     7417 => "00000000",
                     7418 => "00000000",
                     7419 => "00000000",
                     7420 => "00000000",
                     7421 => "00000000",
                     7422 => "00000000",
                     7423 => "00000000",
                     7424 => "00001111",
                     7425 => "00011111",
                     7426 => "00011111",
                     7427 => "00111111",
                     7428 => "00111111",
                     7429 => "01111111",
                     7430 => "01111111",
                     7431 => "01111111",
                     7432 => "11110000",
                     7433 => "11100000",
                     7434 => "11100000",
                     7435 => "11000000",
                     7436 => "11000000",
                     7437 => "10000000",
                     7438 => "10000000",
                     7439 => "10000000",
                     7440 => "11110000",
                     7441 => "11111000",
                     7442 => "11111000",
                     7443 => "11111100",
                     7444 => "11111100",
                     7445 => "11111110",
                     7446 => "11111110",
                     7447 => "11111110",
                     7448 => "00001111",
                     7449 => "00000111",
                     7450 => "00000111",
                     7451 => "00000011",
                     7452 => "00000011",
                     7453 => "00000001",
                     7454 => "00000001",
                     7455 => "00000001",
                     7456 => "01111111",
                     7457 => "01111111",
                     7458 => "00111111",
                     7459 => "00111111",
                     7460 => "00111111",
                     7461 => "00111111",
                     7462 => "00011111",
                     7463 => "00011111",
                     7464 => "10000000",
                     7465 => "10000000",
                     7466 => "11000000",
                     7467 => "11000000",
                     7468 => "11100000",
                     7469 => "11111000",
                     7470 => "11111110",
                     7471 => "11111111",
                     7472 => "11111110",
                     7473 => "11111111",
                     7474 => "11111111",
                     7475 => "11111111",
                     7476 => "11111100",
                     7477 => "11111100",
                     7478 => "11111110",
                     7479 => "11111110",
                     7480 => "11111111",
                     7481 => "01111111",
                     7482 => "00011111",
                     7483 => "00000111",
                     7484 => "00000011",
                     7485 => "00000011",
                     7486 => "00000001",
                     7487 => "10000001",
                     7488 => "01111111",
                     7489 => "01111111",
                     7490 => "01111111",
                     7491 => "00111111",
                     7492 => "00111111",
                     7493 => "00111111",
                     7494 => "00111111",
                     7495 => "00011111",
                     7496 => "10000000",
                     7497 => "10000000",
                     7498 => "10000000",
                     7499 => "11000000",
                     7500 => "11000000",
                     7501 => "11100000",
                     7502 => "11100000",
                     7503 => "11110000",
                     7504 => "11111110",
                     7505 => "11111110",
                     7506 => "11111111",
                     7507 => "11111111",
                     7508 => "11111111",
                     7509 => "11111111",
                     7510 => "11111111",
                     7511 => "11111110",
                     7512 => "00000001",
                     7513 => "00000001",
                     7514 => "00000001",
                     7515 => "00000011",
                     7516 => "00000011",
                     7517 => "00000111",
                     7518 => "00000111",
                     7519 => "00001111",
                     7520 => "00011111",
                     7521 => "00001111",
                     7522 => "00001111",
                     7523 => "00000111",
                     7524 => "00000000",
                     7525 => "00000000",
                     7526 => "00000000",
                     7527 => "00000000",
                     7528 => "11111111",
                     7529 => "11111111",
                     7530 => "11111111",
                     7531 => "11111111",
                     7532 => "11111111",
                     7533 => "11111111",
                     7534 => "11111111",
                     7535 => "11111111",
                     7536 => "11111110",
                     7537 => "11111100",
                     7538 => "11111100",
                     7539 => "11111000",
                     7540 => "00000000",
                     7541 => "00000000",
                     7542 => "00000000",
                     7543 => "00000000",
                     7544 => "11111111",
                     7545 => "11111111",
                     7546 => "11111111",
                     7547 => "11111111",
                     7548 => "11111111",
                     7549 => "11111111",
                     7550 => "11111111",
                     7551 => "11111111",
                     7552 => "01111110",
                     7553 => "01111110",
                     7554 => "01111110",
                     7555 => "01111110",
                     7556 => "01111111",
                     7557 => "01111111",
                     7558 => "01111111",
                     7559 => "01111111",
                     7560 => "10000001",
                     7561 => "10000001",
                     7562 => "10000001",
                     7563 => "10000001",
                     7564 => "10000001",
                     7565 => "10000001",
                     7566 => "10000001",
                     7567 => "10000001",
                     7568 => "11111111",
                     7569 => "11111111",
                     7570 => "11111111",
                     7571 => "11111111",
                     7572 => "11111111",
                     7573 => "11111111",
                     7574 => "11111111",
                     7575 => "11111110",
                     7576 => "00000001",
                     7577 => "00000001",
                     7578 => "00000001",
                     7579 => "00000011",
                     7580 => "00000011",
                     7581 => "00000111",
                     7582 => "00000111",
                     7583 => "00001111",
                     7584 => "11111110",
                     7585 => "11111110",
                     7586 => "11111110",
                     7587 => "11111110",
                     7588 => "11111111",
                     7589 => "11111111",
                     7590 => "11111111",
                     7591 => "11111111",
                     7592 => "00000001",
                     7593 => "00000001",
                     7594 => "00000001",
                     7595 => "00000001",
                     7596 => "00000001",
                     7597 => "00000001",
                     7598 => "00000001",
                     7599 => "00000001",
                     7600 => "01111111",
                     7601 => "01111111",
                     7602 => "01111111",
                     7603 => "01111111",
                     7604 => "01111111",
                     7605 => "01111111",
                     7606 => "01111111",
                     7607 => "01111111",
                     7608 => "10000001",
                     7609 => "10000001",
                     7610 => "10000001",
                     7611 => "10000001",
                     7612 => "10000001",
                     7613 => "10000001",
                     7614 => "10000001",
                     7615 => "10000001",
                     7616 => "11111111",
                     7617 => "11111111",
                     7618 => "11111111",
                     7619 => "11111111",
                     7620 => "11111100",
                     7621 => "11111110",
                     7622 => "11111110",
                     7623 => "01111110",
                     7624 => "11111111",
                     7625 => "00000011",
                     7626 => "00000011",
                     7627 => "00000011",
                     7628 => "00000011",
                     7629 => "00000011",
                     7630 => "00000011",
                     7631 => "11111111",
                     7632 => "11111111",
                     7633 => "11111111",
                     7634 => "11111111",
                     7635 => "11111111",
                     7636 => "00000000",
                     7637 => "00000000",
                     7638 => "00000000",
                     7639 => "00000000",
                     7640 => "11111111",
                     7641 => "11111111",
                     7642 => "11111111",
                     7643 => "11111111",
                     7644 => "11111111",
                     7645 => "11111111",
                     7646 => "11111111",
                     7647 => "11111111",
                     7648 => "01111111",
                     7649 => "01111111",
                     7650 => "01111111",
                     7651 => "01111111",
                     7652 => "01111111",
                     7653 => "01111111",
                     7654 => "01111111",
                     7655 => "01111111",
                     7656 => "10000000",
                     7657 => "10000000",
                     7658 => "10000000",
                     7659 => "10000000",
                     7660 => "10000000",
                     7661 => "10000000",
                     7662 => "10000000",
                     7663 => "10000000",
                     7664 => "11111111",
                     7665 => "11111111",
                     7666 => "11111111",
                     7667 => "11111111",
                     7668 => "11111111",
                     7669 => "11111111",
                     7670 => "11111111",
                     7671 => "11111110",
                     7672 => "00000001",
                     7673 => "00000001",
                     7674 => "00000001",
                     7675 => "00000011",
                     7676 => "00000111",
                     7677 => "00000011",
                     7678 => "00000001",
                     7679 => "00000001",
                     7680 => "01111110",
                     7681 => "01111110",
                     7682 => "01111111",
                     7683 => "01111111",
                     7684 => "01111111",
                     7685 => "01111111",
                     7686 => "01111111",
                     7687 => "01111111",
                     7688 => "10000001",
                     7689 => "10000001",
                     7690 => "10000001",
                     7691 => "10000001",
                     7692 => "10000001",
                     7693 => "10000001",
                     7694 => "10000001",
                     7695 => "10000001",
                     7696 => "00111111",
                     7697 => "00111111",
                     7698 => "00111111",
                     7699 => "00111111",
                     7700 => "00000000",
                     7701 => "00000000",
                     7702 => "00000000",
                     7703 => "00000000",
                     7704 => "11111111",
                     7705 => "11111111",
                     7706 => "11111111",
                     7707 => "11111111",
                     7708 => "11111111",
                     7709 => "11111111",
                     7710 => "11111111",
                     7711 => "11111111",
                     7712 => "01111110",
                     7713 => "01111100",
                     7714 => "01111100",
                     7715 => "01111000",
                     7716 => "00000000",
                     7717 => "00000000",
                     7718 => "00000000",
                     7719 => "00000000",
                     7720 => "11111111",
                     7721 => "11111111",
                     7722 => "11111111",
                     7723 => "11111111",
                     7724 => "11111111",
                     7725 => "11111111",
                     7726 => "11111111",
                     7727 => "11111111",
                     7728 => "11111110",
                     7729 => "11111110",
                     7730 => "11111111",
                     7731 => "11111111",
                     7732 => "01111111",
                     7733 => "01111111",
                     7734 => "01111111",
                     7735 => "01111111",
                     7736 => "10000001",
                     7737 => "10000001",
                     7738 => "10000001",
                     7739 => "10000001",
                     7740 => "10000001",
                     7741 => "10000001",
                     7742 => "10000001",
                     7743 => "10000001",
                     7744 => "01111111",
                     7745 => "01111111",
                     7746 => "00111111",
                     7747 => "00111111",
                     7748 => "00111111",
                     7749 => "00111111",
                     7750 => "00011111",
                     7751 => "00011111",
                     7752 => "10000000",
                     7753 => "10000000",
                     7754 => "11000000",
                     7755 => "11000000",
                     7756 => "11100000",
                     7757 => "11111000",
                     7758 => "11111110",
                     7759 => "11111111",
                     7760 => "00111111",
                     7761 => "10111111",
                     7762 => "11111111",
                     7763 => "11111111",
                     7764 => "11111100",
                     7765 => "11111100",
                     7766 => "11111110",
                     7767 => "11111110",
                     7768 => "11111111",
                     7769 => "01111111",
                     7770 => "00011111",
                     7771 => "00000111",
                     7772 => "00000011",
                     7773 => "00000011",
                     7774 => "00000001",
                     7775 => "10000001",
                     7776 => "01111111",
                     7777 => "01111111",
                     7778 => "01111110",
                     7779 => "01111110",
                     7780 => "01111111",
                     7781 => "01111111",
                     7782 => "01111111",
                     7783 => "01111111",
                     7784 => "10000001",
                     7785 => "10000001",
                     7786 => "10000001",
                     7787 => "10000001",
                     7788 => "10000001",
                     7789 => "10000001",
                     7790 => "10000001",
                     7791 => "10000001",
                     7792 => "01111110",
                     7793 => "01111110",
                     7794 => "01111110",
                     7795 => "01111110",
                     7796 => "01111111",
                     7797 => "01111111",
                     7798 => "01111111",
                     7799 => "01111111",
                     7800 => "10000001",
                     7801 => "10000001",
                     7802 => "10000001",
                     7803 => "10000001",
                     7804 => "10000001",
                     7805 => "10000001",
                     7806 => "10000001",
                     7807 => "10000001",
                     7808 => "10000001",
                     7809 => "11000011",
                     7810 => "11000011",
                     7811 => "11100111",
                     7812 => "11100111",
                     7813 => "11111111",
                     7814 => "11111111",
                     7815 => "11111111",
                     7816 => "01111110",
                     7817 => "00111100",
                     7818 => "00111100",
                     7819 => "00011000",
                     7820 => "00011000",
                     7821 => "00000000",
                     7822 => "00000000",
                     7823 => "00000000",
                     7824 => "00001111",
                     7825 => "01000011",
                     7826 => "01011011",
                     7827 => "01010011",
                     7828 => "00110001",
                     7829 => "00011001",
                     7830 => "00001111",
                     7831 => "00000111",
                     7832 => "11110010",
                     7833 => "11111110",
                     7834 => "11111110",
                     7835 => "11111111",
                     7836 => "11111111",
                     7837 => "11101111",
                     7838 => "11110111",
                     7839 => "11111000",
                     7840 => "11000001",
                     7841 => "11000011",
                     7842 => "11000110",
                     7843 => "10000100",
                     7844 => "11111100",
                     7845 => "11111100",
                     7846 => "00001110",
                     7847 => "00000010",
                     7848 => "10111111",
                     7849 => "10111110",
                     7850 => "10111101",
                     7851 => "01111011",
                     7852 => "01111011",
                     7853 => "00000111",
                     7854 => "11110011",
                     7855 => "11111101",
                     7856 => "00010000",
                     7857 => "00100000",
                     7858 => "00100010",
                     7859 => "10111010",
                     7860 => "11100110",
                     7861 => "11100001",
                     7862 => "11000000",
                     7863 => "11000000",
                     7864 => "11111111",
                     7865 => "11111111",
                     7866 => "11111111",
                     7867 => "01100111",
                     7868 => "01011001",
                     7869 => "10011110",
                     7870 => "10111111",
                     7871 => "10111111",
                     7872 => "00100000",
                     7873 => "10100110",
                     7874 => "01010100",
                     7875 => "00100110",
                     7876 => "00100000",
                     7877 => "11000110",
                     7878 => "01010100",
                     7879 => "00100110",
                     7880 => "00100000",
                     7881 => "11100110",
                     7882 => "01010100",
                     7883 => "00100110",
                     7884 => "00100001",
                     7885 => "00000110",
                     7886 => "01010100",
                     7887 => "00100110",
                     7888 => "00100000",
                     7889 => "10000101",
                     7890 => "00000001",
                     7891 => "01000100",
                     7892 => "00100000",
                     7893 => "10000110",
                     7894 => "01010100",
                     7895 => "01001000",
                     7896 => "00100000",
                     7897 => "10011010",
                     7898 => "00000001",
                     7899 => "01001001",
                     7900 => "00100000",
                     7901 => "10100101",
                     7902 => "11001001",
                     7903 => "01000110",
                     7904 => "00100000",
                     7905 => "10111010",
                     7906 => "11001001",
                     7907 => "01001010",
                     7908 => "00100000",
                     7909 => "10100110",
                     7910 => "00001010",
                     7911 => "11010000",
                     7912 => "11010001",
                     7913 => "11011000",
                     7914 => "11011000",
                     7915 => "11011110",
                     7916 => "11010001",
                     7917 => "11010000",
                     7918 => "11011010",
                     7919 => "11011110",
                     7920 => "11010001",
                     7921 => "00100000",
                     7922 => "11000110",
                     7923 => "00001010",
                     7924 => "11010010",
                     7925 => "11010011",
                     7926 => "11011011",
                     7927 => "11011011",
                     7928 => "11011011",
                     7929 => "11011001",
                     7930 => "11011011",
                     7931 => "11011100",
                     7932 => "11011011",
                     7933 => "11011111",
                     7934 => "00100000",
                     7935 => "11100110",
                     7936 => "00001010",
                     7937 => "11010100",
                     7938 => "11010101",
                     7939 => "11010100",
                     7940 => "11011001",
                     7941 => "11011011",
                     7942 => "11100010",
                     7943 => "11010100",
                     7944 => "11011010",
                     7945 => "11011011",
                     7946 => "11100000",
                     7947 => "00100001",
                     7948 => "00000110",
                     7949 => "00001010",
                     7950 => "11010110",
                     7951 => "11010111",
                     7952 => "11010110",
                     7953 => "11010111",
                     7954 => "11100001",
                     7955 => "00100110",
                     7956 => "11010110",
                     7957 => "11011101",
                     7958 => "11100001",
                     7959 => "11100001",
                     7960 => "00100001",
                     7961 => "00100110",
                     7962 => "00010100",
                     7963 => "11010000",
                     7964 => "11101000",
                     7965 => "11010001",
                     7966 => "11010000",
                     7967 => "11010001",
                     7968 => "11011110",
                     7969 => "11010001",
                     7970 => "11011000",
                     7971 => "11010000",
                     7972 => "11010001",
                     7973 => "00100110",
                     7974 => "11011110",
                     7975 => "11010001",
                     7976 => "11011110",
                     7977 => "11010001",
                     7978 => "11010000",
                     7979 => "11010001",
                     7980 => "11010000",
                     7981 => "11010001",
                     7982 => "00100110",
                     7983 => "00100001",
                     7984 => "01000110",
                     7985 => "00010100",
                     7986 => "11011011",
                     7987 => "01000010",
                     7988 => "01000010",
                     7989 => "11011011",
                     7990 => "01000010",
                     7991 => "11011011",
                     7992 => "01000010",
                     7993 => "11011011",
                     7994 => "11011011",
                     7995 => "01000010",
                     7996 => "00100110",
                     7997 => "11011011",
                     7998 => "01000010",
                     7999 => "11011011",
                     8000 => "01000010",
                     8001 => "11011011",
                     8002 => "01000010",
                     8003 => "11011011",
                     8004 => "01000010",
                     8005 => "00100110",
                     8006 => "00100001",
                     8007 => "01100110",
                     8008 => "01000110",
                     8009 => "11011011",
                     8010 => "00100001",
                     8011 => "01101100",
                     8012 => "00001110",
                     8013 => "11011111",
                     8014 => "11011011",
                     8015 => "11011011",
                     8016 => "11011011",
                     8017 => "00100110",
                     8018 => "11011011",
                     8019 => "11011111",
                     8020 => "11011011",
                     8021 => "11011111",
                     8022 => "11011011",
                     8023 => "11011011",
                     8024 => "11100100",
                     8025 => "11100101",
                     8026 => "00100110",
                     8027 => "00100001",
                     8028 => "10000110",
                     8029 => "00010100",
                     8030 => "11011011",
                     8031 => "11011011",
                     8032 => "11011011",
                     8033 => "11011110",
                     8034 => "01000011",
                     8035 => "11011011",
                     8036 => "11100000",
                     8037 => "11011011",
                     8038 => "11011011",
                     8039 => "11011011",
                     8040 => "00100110",
                     8041 => "11011011",
                     8042 => "11100011",
                     8043 => "11011011",
                     8044 => "11100000",
                     8045 => "11011011",
                     8046 => "11011011",
                     8047 => "11100110",
                     8048 => "11100011",
                     8049 => "00100110",
                     8050 => "00100001",
                     8051 => "10100110",
                     8052 => "00010100",
                     8053 => "11011011",
                     8054 => "11011011",
                     8055 => "11011011",
                     8056 => "11011011",
                     8057 => "01000010",
                     8058 => "11011011",
                     8059 => "11011011",
                     8060 => "11011011",
                     8061 => "11010100",
                     8062 => "11011001",
                     8063 => "00100110",
                     8064 => "11011011",
                     8065 => "11011001",
                     8066 => "11011011",
                     8067 => "11011011",
                     8068 => "11010100",
                     8069 => "11011001",
                     8070 => "11010100",
                     8071 => "11011001",
                     8072 => "11100111",
                     8073 => "00100001",
                     8074 => "11000101",
                     8075 => "00010110",
                     8076 => "01011111",
                     8077 => "10010101",
                     8078 => "10010101",
                     8079 => "10010101",
                     8080 => "10010101",
                     8081 => "10010101",
                     8082 => "10010101",
                     8083 => "10010101",
                     8084 => "10010101",
                     8085 => "10010111",
                     8086 => "10011000",
                     8087 => "01111000",
                     8088 => "10010101",
                     8089 => "10010110",
                     8090 => "10010101",
                     8091 => "10010101",
                     8092 => "10010111",
                     8093 => "10011000",
                     8094 => "10010111",
                     8095 => "10011000",
                     8096 => "10010101",
                     8097 => "01111010",
                     8098 => "00100001",
                     8099 => "11101101",
                     8100 => "00001110",
                     8101 => "11001111",
                     8102 => "00000001",
                     8103 => "00001001",
                     8104 => "00001000",
                     8105 => "00000101",
                     8106 => "00100100",
                     8107 => "00010111",
                     8108 => "00010010",
                     8109 => "00010111",
                     8110 => "00011101",
                     8111 => "00001110",
                     8112 => "00010111",
                     8113 => "00001101",
                     8114 => "00011000",
                     8115 => "00100010",
                     8116 => "01001011",
                     8117 => "00001101",
                     8118 => "00000001",
                     8119 => "00100100",
                     8120 => "00011001",
                     8121 => "00010101",
                     8122 => "00001010",
                     8123 => "00100010",
                     8124 => "00001110",
                     8125 => "00011011",
                     8126 => "00100100",
                     8127 => "00010000",
                     8128 => "00001010",
                     8129 => "00010110",
                     8130 => "00001110",
                     8131 => "00100010",
                     8132 => "10001011",
                     8133 => "00001101",
                     8134 => "00000010",
                     8135 => "00100100",
                     8136 => "00011001",
                     8137 => "00010101",
                     8138 => "00001010",
                     8139 => "00100010",
                     8140 => "00001110",
                     8141 => "00011011",
                     8142 => "00100100",
                     8143 => "00010000",
                     8144 => "00001010",
                     8145 => "00010110",
                     8146 => "00001110",
                     8147 => "00100010",
                     8148 => "11101100",
                     8149 => "00000100",
                     8150 => "00011101",
                     8151 => "00011000",
                     8152 => "00011001",
                     8153 => "00101000",
                     8154 => "00100010",
                     8155 => "11110110",
                     8156 => "00000001",
                     8157 => "00000000",
                     8158 => "00100011",
                     8159 => "11001001",
                     8160 => "01010110",
                     8161 => "01010101",
                     8162 => "00100011",
                     8163 => "11100010",
                     8164 => "00000100",
                     8165 => "10011001",
                     8166 => "10101010",
                     8167 => "10101010",
                     8168 => "10101010",
                     8169 => "00100011",
                     8170 => "11101010",
                     8171 => "00000100",
                     8172 => "10011001",
                     8173 => "10101010",
                     8174 => "10101010",
                     8175 => "10101010",
                     8176 => "00000000",
                     8177 => "11111111",
                     8178 => "11111111",
                     8179 => "11111111",
                     8180 => "11111111",
                     8181 => "11111111",
                     8182 => "11111111",
                     8183 => "11111111",
                     8184 => "11111111",
                     8185 => "11111111",
                     8186 => "11111111",
                     8187 => "11111111",
                     8188 => "11111111",
                     8189 => "11111111",
                     8190 => "11111111",
                     8191 => "11111111"
                    );
            else
                --ProgramData <= prg_rom(conv_integer(to_unsigned(ProgramAddress, ProgramAddress'length)));
                --CharacterData <= chr_rom(conv_integer(to_unsigned(CharacterAddress, CharacterAddress'length)));
            end if;
				
				
				ProgramData <= prg_rom(to_integer(unsigned(ProgramAddress)));
				CharacterData <= chr_rom(to_integer(unsigned(CharacterAddress)));
        end if;
    end process;

end arch;

